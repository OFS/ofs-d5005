// Copyright 2021 Intel Corporation
// SPDX-License-Identifier: MIT

//-----------------------------------------------------------------------------
// Description : Contains all sequences 
//-----------------------------------------------------------------------------

`ifndef SEQ_LIB_SVH
`define SEQ_LIB_SVH

`include "pcie_hip_defines.svh"
`include "pcie_device_report_catcher.sv"
`include "vip_seq/enumerate_seq.sv"
`include "pcie_vip_seq.svh"
`include "pcie_device_sequence_library.sv"
`include "vip_seq/flr_rst_seq.sv"
`include "axi_slave_mem_response_sequence.sv"
`include "axi_simple_reset_sequence.sv"
`include "config_seq.svh"
`include "base_seq.svh"
`include "mmio_seq.svh"
`include "he_lpbk_seq.svh"
`include "he_lpbk_long_seq.svh"
`include "he_lpbk_rd_seq.svh"
`include "he_lpbk_wr_seq.svh"
`include "he_lpbk_thruput_seq.svh"
`include "he_lpbk_rd_cont_seq.svh"
`include "he_lpbk_wr_cont_seq.svh"
`include "he_lpbk_thruput_contmode_seq.svh"
`include "he_mem_lpbk_seq.svh"
`include "he_mem_lpbk_long_seq.svh"
`include "he_mem_rd_seq.svh"
`include "he_mem_wr_seq.svh"
`include "he_mem_thruput_seq.svh"
`include "he_mem_rd_cont_seq.svh"
`include "he_mem_wr_cont_seq.svh"
`include "he_mem_thruput_contmode_seq.svh"
`include "he_mem_cont_seq.svh"
`include "he_hssi_tx_lpbk.svh"
`include "he_hssi_err_seq.svh"
`include "he_hssi_csr_seq.svh"
`include "mmio_stress_seq.svh"
`include "he_random_seq.svh"
`include "dfh_walking_seq.svh"
`include "mmio_unimp_seq.svh"
`include "he_lpbk_reqlen1_seq.svh"
`include "he_lpbk_reqlen2_seq.svh"
`include "he_lpbk_reqlen4_seq.svh"
`include "he_lpbk_reqlen8_seq.svh"
`include "he_mem_lpbk_reqlen1_seq.svh"
`include "he_mem_lpbk_reqlen2_seq.svh"
`include "he_mem_lpbk_reqlen4_seq.svh"
`include "he_lpbk_long_rst_seq.svh"
`include "he_mem_lpbk_long_rst_seq.svh"
`include "mmio_stress_nonblocking_seq.svh"
`include "he_lpbk_cont_seq.svh"
`include "fme_csr_seq.svh"
`include "msix_csr_seq.svh"
`include "pmci_csr_seq.svh"
`include "helb_csr_seq.svh"
`include "hemem_csr_seq.svh"
`include "hehssi_csr_seq.svh"
`include "mini_smoke_seq.svh"
`include "fme_intr_seq.svh"
`include "flr_reset_seq.svh"
`include "flr_vf0_reset_seq.svh"
`include "flr_vf1_reset_seq.svh"
`include "flr_vf2_reset_seq.svh"
`include "port_gasket_csr_seq.svh"
`include "helb_rd_1cl_seq.svh"
`include "helb_rd_2cl_seq.svh"
`include "helb_rd_4cl_seq.svh"
`include "helb_wr_1cl_seq.svh"
`include "helb_wr_2cl_seq.svh"
`include "helb_wr_4cl_seq.svh"
`include "helb_thruput_1cl_seq.svh"
`include "helb_thruput_2cl_seq.svh"
`include "helb_thruput_4cl_seq.svh"
`include "he_random_long_seq.svh"
`include "hemem_intr_seq.svh"
`include "he_lpbk_port_rst_seq.svh"
`include "he_hssi_rx_lpbk.svh"
`include "fme_ras_cat_fat_err_seq.svh"
`include "fme_ras_no_fat_err_seq.svh"
`include "protocol_checker_csr_seq.svh"
`include "MaxTagError_seq.svh"
`include "TxMWrDataPayloadOverrun_seq.svh"
`include "TxMWrInsufficientData_seq.svh"
`include "UnexpMMIORspErr_seq.svh"
`include "malformedtlp_seq.svh"
`include "maxpayloaderror_seq.svh"
`include "MMIOInsufficientData_seq.svh"
`include "MMIOTimedOut_seq.svh"
`include "MMIODataPayloadOverrun_seq.svh"
`include "he_user_intr_seq.svh"
`include "he_mem_user_intr_seq.svh"
`include "he_mem_multi_user_intr_seq.svh"

`endif // SEQ_LIB_SVH
