// Copyright 2020 Intel Corporation
// SPDX-License-Identifier: MIT

// DUT_pcie_tb_ip.v

// Generated using ACDS version 19.2 57

`timescale 1 ps / 1 ps
module DUT_pcie_tb_ip #(
		parameter lane_mask_hwtcl                      = "x16",
		parameter pll_refclk_freq_hwtcl                = "100 MHz",
		parameter serial_sim_hwtcl                     = 1,
		parameter deemphasis_enable_hwtcl              = "false",
		parameter pld_clk_MHz                          = 125,
		parameter millisecond_cycle_count_hwtcl        = 124250,
		parameter use_crc_forwarding_hwtcl             = 0,
		parameter ecrc_check_capable_hwtcl             = 0,
		parameter ecrc_gen_capable_hwtcl               = 0,
		parameter bfm_drive_interface_clk_hwtcl        = 1,
		parameter bfm_drive_interface_npor_hwtcl       = 1,
		parameter bfm_drive_interface_pipe_hwtcl       = 1,
		parameter bfm_drive_interface_control_hwtcl    = 1,
		parameter select_example_design_sim_BFM_hwtcl  = "Intel FPGA BFM",
		parameter enable_pipe32_phyip_ser_driver_hwtcl = 0
	) (
		output wire        rx_in0,                    // hip_serial.rx_in0
		output wire        rx_in1,                    //           .rx_in1
		output wire        rx_in2,                    //           .rx_in2
		output wire        rx_in3,                    //           .rx_in3
		output wire        rx_in4,                    //           .rx_in4
		output wire        rx_in5,                    //           .rx_in5
		output wire        rx_in6,                    //           .rx_in6
		output wire        rx_in7,                    //           .rx_in7
		output wire        rx_in8,                    //           .rx_in8
		output wire        rx_in9,                    //           .rx_in9
		output wire        rx_in10,                   //           .rx_in10
		output wire        rx_in11,                   //           .rx_in11
		output wire        rx_in12,                   //           .rx_in12
		output wire        rx_in13,                   //           .rx_in13
		output wire        rx_in14,                   //           .rx_in14
		output wire        rx_in15,                   //           .rx_in15
		input  wire        tx_out0,                   //           .tx_out0
		input  wire        tx_out1,                   //           .tx_out1
		input  wire        tx_out2,                   //           .tx_out2
		input  wire        tx_out3,                   //           .tx_out3
		input  wire        tx_out4,                   //           .tx_out4
		input  wire        tx_out5,                   //           .tx_out5
		input  wire        tx_out6,                   //           .tx_out6
		input  wire        tx_out7,                   //           .tx_out7
		input  wire        tx_out8,                   //           .tx_out8
		input  wire        tx_out9,                   //           .tx_out9
		input  wire        tx_out10,                  //           .tx_out10
		input  wire        tx_out11,                  //           .tx_out11
		input  wire        tx_out12,                  //           .tx_out12
		input  wire        tx_out13,                  //           .tx_out13
		input  wire        tx_out14,                  //           .tx_out14
		input  wire        tx_out15,                  //           .tx_out15
		output wire        refclk,                    //     refclk.clk
		output wire        sim_pipe_pclk_in,          //   hip_pipe.sim_pipe_pclk_in
		output wire        sim_pipe_mask_tx_pll_lock, //           .sim_pipe_mask_tx_pll_lock
		input  wire [1:0]  sim_pipe_rate,             //           .sim_pipe_rate
		input  wire [5:0]  sim_ltssmstate,            //           .sim_ltssmstate
		output wire [5:0]  dirfeedback0,              //           .dirfeedback0
		output wire [5:0]  dirfeedback1,              //           .dirfeedback1
		output wire [5:0]  dirfeedback2,              //           .dirfeedback2
		output wire [5:0]  dirfeedback3,              //           .dirfeedback3
		output wire [5:0]  dirfeedback4,              //           .dirfeedback4
		output wire [5:0]  dirfeedback5,              //           .dirfeedback5
		output wire [5:0]  dirfeedback6,              //           .dirfeedback6
		output wire [5:0]  dirfeedback7,              //           .dirfeedback7
		input  wire        rxeqeval0,                 //           .rxeqeval0
		input  wire        rxeqeval1,                 //           .rxeqeval1
		input  wire        rxeqeval2,                 //           .rxeqeval2
		input  wire        rxeqeval3,                 //           .rxeqeval3
		input  wire        rxeqeval4,                 //           .rxeqeval4
		input  wire        rxeqeval5,                 //           .rxeqeval5
		input  wire        rxeqeval6,                 //           .rxeqeval6
		input  wire        rxeqeval7,                 //           .rxeqeval7
		input  wire        rxeqinprogress0,           //           .rxeqinprogress0
		input  wire        rxeqinprogress1,           //           .rxeqinprogress1
		input  wire        rxeqinprogress2,           //           .rxeqinprogress2
		input  wire        rxeqinprogress3,           //           .rxeqinprogress3
		input  wire        rxeqinprogress4,           //           .rxeqinprogress4
		input  wire        rxeqinprogress5,           //           .rxeqinprogress5
		input  wire        rxeqinprogress6,           //           .rxeqinprogress6
		input  wire        rxeqinprogress7,           //           .rxeqinprogress7
		input  wire        invalidreq0,               //           .invalidreq0
		input  wire        invalidreq1,               //           .invalidreq1
		input  wire        invalidreq2,               //           .invalidreq2
		input  wire        invalidreq3,               //           .invalidreq3
		input  wire        invalidreq4,               //           .invalidreq4
		input  wire        invalidreq5,               //           .invalidreq5
		input  wire        invalidreq6,               //           .invalidreq6
		input  wire        invalidreq7,               //           .invalidreq7
		input  wire [1:0]  powerdown0,                //           .powerdown0
		input  wire [1:0]  powerdown1,                //           .powerdown1
		input  wire [1:0]  powerdown2,                //           .powerdown2
		input  wire [1:0]  powerdown3,                //           .powerdown3
		input  wire [1:0]  powerdown4,                //           .powerdown4
		input  wire [1:0]  powerdown5,                //           .powerdown5
		input  wire [1:0]  powerdown6,                //           .powerdown6
		input  wire [1:0]  powerdown7,                //           .powerdown7
		input  wire        rxpolarity0,               //           .rxpolarity0
		input  wire        rxpolarity1,               //           .rxpolarity1
		input  wire        rxpolarity2,               //           .rxpolarity2
		input  wire        rxpolarity3,               //           .rxpolarity3
		input  wire        rxpolarity4,               //           .rxpolarity4
		input  wire        rxpolarity5,               //           .rxpolarity5
		input  wire        rxpolarity6,               //           .rxpolarity6
		input  wire        rxpolarity7,               //           .rxpolarity7
		input  wire        txcompl0,                  //           .txcompl0
		input  wire        txcompl1,                  //           .txcompl1
		input  wire        txcompl2,                  //           .txcompl2
		input  wire        txcompl3,                  //           .txcompl3
		input  wire        txcompl4,                  //           .txcompl4
		input  wire        txcompl5,                  //           .txcompl5
		input  wire        txcompl6,                  //           .txcompl6
		input  wire        txcompl7,                  //           .txcompl7
		input  wire [31:0] txdata0,                   //           .txdata0
		input  wire [31:0] txdata1,                   //           .txdata1
		input  wire [31:0] txdata2,                   //           .txdata2
		input  wire [31:0] txdata3,                   //           .txdata3
		input  wire [31:0] txdata4,                   //           .txdata4
		input  wire [31:0] txdata5,                   //           .txdata5
		input  wire [31:0] txdata6,                   //           .txdata6
		input  wire [31:0] txdata7,                   //           .txdata7
		input  wire [3:0]  txdatak0,                  //           .txdatak0
		input  wire [3:0]  txdatak1,                  //           .txdatak1
		input  wire [3:0]  txdatak2,                  //           .txdatak2
		input  wire [3:0]  txdatak3,                  //           .txdatak3
		input  wire [3:0]  txdatak4,                  //           .txdatak4
		input  wire [3:0]  txdatak5,                  //           .txdatak5
		input  wire [3:0]  txdatak6,                  //           .txdatak6
		input  wire [3:0]  txdatak7,                  //           .txdatak7
		input  wire        txdetectrx0,               //           .txdetectrx0
		input  wire        txdetectrx1,               //           .txdetectrx1
		input  wire        txdetectrx2,               //           .txdetectrx2
		input  wire        txdetectrx3,               //           .txdetectrx3
		input  wire        txdetectrx4,               //           .txdetectrx4
		input  wire        txdetectrx5,               //           .txdetectrx5
		input  wire        txdetectrx6,               //           .txdetectrx6
		input  wire        txdetectrx7,               //           .txdetectrx7
		input  wire        txelecidle0,               //           .txelecidle0
		input  wire        txelecidle1,               //           .txelecidle1
		input  wire        txelecidle2,               //           .txelecidle2
		input  wire        txelecidle3,               //           .txelecidle3
		input  wire        txelecidle4,               //           .txelecidle4
		input  wire        txelecidle5,               //           .txelecidle5
		input  wire        txelecidle6,               //           .txelecidle6
		input  wire        txelecidle7,               //           .txelecidle7
		input  wire        txdeemph0,                 //           .txdeemph0
		input  wire        txdeemph1,                 //           .txdeemph1
		input  wire        txdeemph2,                 //           .txdeemph2
		input  wire        txdeemph3,                 //           .txdeemph3
		input  wire        txdeemph4,                 //           .txdeemph4
		input  wire        txdeemph5,                 //           .txdeemph5
		input  wire        txdeemph6,                 //           .txdeemph6
		input  wire        txdeemph7,                 //           .txdeemph7
		input  wire [2:0]  txmargin0,                 //           .txmargin0
		input  wire [2:0]  txmargin1,                 //           .txmargin1
		input  wire [2:0]  txmargin2,                 //           .txmargin2
		input  wire [2:0]  txmargin3,                 //           .txmargin3
		input  wire [2:0]  txmargin4,                 //           .txmargin4
		input  wire [2:0]  txmargin5,                 //           .txmargin5
		input  wire [2:0]  txmargin6,                 //           .txmargin6
		input  wire [2:0]  txmargin7,                 //           .txmargin7
		input  wire        txswing0,                  //           .txswing0
		input  wire        txswing1,                  //           .txswing1
		input  wire        txswing2,                  //           .txswing2
		input  wire        txswing3,                  //           .txswing3
		input  wire        txswing4,                  //           .txswing4
		input  wire        txswing5,                  //           .txswing5
		input  wire        txswing6,                  //           .txswing6
		input  wire        txswing7,                  //           .txswing7
		output wire        phystatus0,                //           .phystatus0
		output wire        phystatus1,                //           .phystatus1
		output wire        phystatus2,                //           .phystatus2
		output wire        phystatus3,                //           .phystatus3
		output wire        phystatus4,                //           .phystatus4
		output wire        phystatus5,                //           .phystatus5
		output wire        phystatus6,                //           .phystatus6
		output wire        phystatus7,                //           .phystatus7
		output wire [31:0] rxdata0,                   //           .rxdata0
		output wire [31:0] rxdata1,                   //           .rxdata1
		output wire [31:0] rxdata2,                   //           .rxdata2
		output wire [31:0] rxdata3,                   //           .rxdata3
		output wire [31:0] rxdata4,                   //           .rxdata4
		output wire [31:0] rxdata5,                   //           .rxdata5
		output wire [31:0] rxdata6,                   //           .rxdata6
		output wire [31:0] rxdata7,                   //           .rxdata7
		output wire [3:0]  rxdatak0,                  //           .rxdatak0
		output wire [3:0]  rxdatak1,                  //           .rxdatak1
		output wire [3:0]  rxdatak2,                  //           .rxdatak2
		output wire [3:0]  rxdatak3,                  //           .rxdatak3
		output wire [3:0]  rxdatak4,                  //           .rxdatak4
		output wire [3:0]  rxdatak5,                  //           .rxdatak5
		output wire [3:0]  rxdatak6,                  //           .rxdatak6
		output wire [3:0]  rxdatak7,                  //           .rxdatak7
		output wire        rxelecidle0,               //           .rxelecidle0
		output wire        rxelecidle1,               //           .rxelecidle1
		output wire        rxelecidle2,               //           .rxelecidle2
		output wire        rxelecidle3,               //           .rxelecidle3
		output wire        rxelecidle4,               //           .rxelecidle4
		output wire        rxelecidle5,               //           .rxelecidle5
		output wire        rxelecidle6,               //           .rxelecidle6
		output wire        rxelecidle7,               //           .rxelecidle7
		output wire [2:0]  rxstatus0,                 //           .rxstatus0
		output wire [2:0]  rxstatus1,                 //           .rxstatus1
		output wire [2:0]  rxstatus2,                 //           .rxstatus2
		output wire [2:0]  rxstatus3,                 //           .rxstatus3
		output wire [2:0]  rxstatus4,                 //           .rxstatus4
		output wire [2:0]  rxstatus5,                 //           .rxstatus5
		output wire [2:0]  rxstatus6,                 //           .rxstatus6
		output wire [2:0]  rxstatus7,                 //           .rxstatus7
		output wire        rxvalid0,                  //           .rxvalid0
		output wire        rxvalid1,                  //           .rxvalid1
		output wire        rxvalid2,                  //           .rxvalid2
		output wire        rxvalid3,                  //           .rxvalid3
		output wire        rxvalid4,                  //           .rxvalid4
		output wire        rxvalid5,                  //           .rxvalid5
		output wire        rxvalid6,                  //           .rxvalid6
		output wire        rxvalid7,                  //           .rxvalid7
		output wire        rxdataskip0,               //           .rxdataskip0
		output wire        rxdataskip1,               //           .rxdataskip1
		output wire        rxdataskip2,               //           .rxdataskip2
		output wire        rxdataskip3,               //           .rxdataskip3
		output wire        rxdataskip4,               //           .rxdataskip4
		output wire        rxdataskip5,               //           .rxdataskip5
		output wire        rxdataskip6,               //           .rxdataskip6
		output wire        rxdataskip7,               //           .rxdataskip7
		output wire        rxblkst0,                  //           .rxblkst0
		output wire        rxblkst1,                  //           .rxblkst1
		output wire        rxblkst2,                  //           .rxblkst2
		output wire        rxblkst3,                  //           .rxblkst3
		output wire        rxblkst4,                  //           .rxblkst4
		output wire        rxblkst5,                  //           .rxblkst5
		output wire        rxblkst6,                  //           .rxblkst6
		output wire        rxblkst7,                  //           .rxblkst7
		output wire [1:0]  rxsynchd0,                 //           .rxsynchd0
		output wire [1:0]  rxsynchd1,                 //           .rxsynchd1
		output wire [1:0]  rxsynchd2,                 //           .rxsynchd2
		output wire [1:0]  rxsynchd3,                 //           .rxsynchd3
		output wire [1:0]  rxsynchd4,                 //           .rxsynchd4
		output wire [1:0]  rxsynchd5,                 //           .rxsynchd5
		output wire [1:0]  rxsynchd6,                 //           .rxsynchd6
		output wire [1:0]  rxsynchd7,                 //           .rxsynchd7
		input  wire [17:0] currentcoeff0,             //           .currentcoeff0
		input  wire [17:0] currentcoeff1,             //           .currentcoeff1
		input  wire [17:0] currentcoeff2,             //           .currentcoeff2
		input  wire [17:0] currentcoeff3,             //           .currentcoeff3
		input  wire [17:0] currentcoeff4,             //           .currentcoeff4
		input  wire [17:0] currentcoeff5,             //           .currentcoeff5
		input  wire [17:0] currentcoeff6,             //           .currentcoeff6
		input  wire [17:0] currentcoeff7,             //           .currentcoeff7
		input  wire [2:0]  currentrxpreset0,          //           .currentrxpreset0
		input  wire [2:0]  currentrxpreset1,          //           .currentrxpreset1
		input  wire [2:0]  currentrxpreset2,          //           .currentrxpreset2
		input  wire [2:0]  currentrxpreset3,          //           .currentrxpreset3
		input  wire [2:0]  currentrxpreset4,          //           .currentrxpreset4
		input  wire [2:0]  currentrxpreset5,          //           .currentrxpreset5
		input  wire [2:0]  currentrxpreset6,          //           .currentrxpreset6
		input  wire [2:0]  currentrxpreset7,          //           .currentrxpreset7
		input  wire [1:0]  txsynchd0,                 //           .txsynchd0
		input  wire [1:0]  txsynchd1,                 //           .txsynchd1
		input  wire [1:0]  txsynchd2,                 //           .txsynchd2
		input  wire [1:0]  txsynchd3,                 //           .txsynchd3
		input  wire [1:0]  txsynchd4,                 //           .txsynchd4
		input  wire [1:0]  txsynchd5,                 //           .txsynchd5
		input  wire [1:0]  txsynchd6,                 //           .txsynchd6
		input  wire [1:0]  txsynchd7,                 //           .txsynchd7
		input  wire        txblkst0,                  //           .txblkst0
		input  wire        txblkst1,                  //           .txblkst1
		input  wire        txblkst2,                  //           .txblkst2
		input  wire        txblkst3,                  //           .txblkst3
		input  wire        txblkst4,                  //           .txblkst4
		input  wire        txblkst5,                  //           .txblkst5
		input  wire        txblkst6,                  //           .txblkst6
		input  wire        txblkst7,                  //           .txblkst7
		input  wire        txdataskip0,               //           .txdataskip0
		input  wire        txdataskip1,               //           .txdataskip1
		input  wire        txdataskip2,               //           .txdataskip2
		input  wire        txdataskip3,               //           .txdataskip3
		input  wire        txdataskip4,               //           .txdataskip4
		input  wire        txdataskip5,               //           .txdataskip5
		input  wire        txdataskip6,               //           .txdataskip6
		input  wire        txdataskip7,               //           .txdataskip7
		input  wire [1:0]  rate0,                     //           .rate0
		input  wire [1:0]  rate1,                     //           .rate1
		input  wire [1:0]  rate2,                     //           .rate2
		input  wire [1:0]  rate3,                     //           .rate3
		input  wire [1:0]  rate4,                     //           .rate4
		input  wire [1:0]  rate5,                     //           .rate5
		input  wire [1:0]  rate6,                     //           .rate6
		input  wire [1:0]  rate7,                     //           .rate7
		output wire [5:0]  dirfeedback8,              //           .dirfeedback8
		output wire [5:0]  dirfeedback9,              //           .dirfeedback9
		output wire [5:0]  dirfeedback10,             //           .dirfeedback10
		output wire [5:0]  dirfeedback11,             //           .dirfeedback11
		output wire [5:0]  dirfeedback12,             //           .dirfeedback12
		output wire [5:0]  dirfeedback13,             //           .dirfeedback13
		output wire [5:0]  dirfeedback14,             //           .dirfeedback14
		output wire [5:0]  dirfeedback15,             //           .dirfeedback15
		input  wire        rxeqeval8,                 //           .rxeqeval8
		input  wire        rxeqeval9,                 //           .rxeqeval9
		input  wire        rxeqeval10,                //           .rxeqeval10
		input  wire        rxeqeval11,                //           .rxeqeval11
		input  wire        rxeqeval12,                //           .rxeqeval12
		input  wire        rxeqeval13,                //           .rxeqeval13
		input  wire        rxeqeval14,                //           .rxeqeval14
		input  wire        rxeqeval15,                //           .rxeqeval15
		input  wire        rxeqinprogress8,           //           .rxeqinprogress8
		input  wire        rxeqinprogress9,           //           .rxeqinprogress9
		input  wire        rxeqinprogress10,          //           .rxeqinprogress10
		input  wire        rxeqinprogress11,          //           .rxeqinprogress11
		input  wire        rxeqinprogress12,          //           .rxeqinprogress12
		input  wire        rxeqinprogress13,          //           .rxeqinprogress13
		input  wire        rxeqinprogress14,          //           .rxeqinprogress14
		input  wire        rxeqinprogress15,          //           .rxeqinprogress15
		input  wire        invalidreq8,               //           .invalidreq8
		input  wire        invalidreq9,               //           .invalidreq9
		input  wire        invalidreq10,              //           .invalidreq10
		input  wire        invalidreq11,              //           .invalidreq11
		input  wire        invalidreq12,              //           .invalidreq12
		input  wire        invalidreq13,              //           .invalidreq13
		input  wire        invalidreq14,              //           .invalidreq14
		input  wire        invalidreq15,              //           .invalidreq15
		input  wire [1:0]  powerdown8,                //           .powerdown8
		input  wire [1:0]  powerdown9,                //           .powerdown9
		input  wire [1:0]  powerdown10,               //           .powerdown10
		input  wire [1:0]  powerdown11,               //           .powerdown11
		input  wire [1:0]  powerdown12,               //           .powerdown12
		input  wire [1:0]  powerdown13,               //           .powerdown13
		input  wire [1:0]  powerdown14,               //           .powerdown14
		input  wire [1:0]  powerdown15,               //           .powerdown15
		input  wire        rxpolarity8,               //           .rxpolarity8
		input  wire        rxpolarity9,               //           .rxpolarity9
		input  wire        rxpolarity10,              //           .rxpolarity10
		input  wire        rxpolarity11,              //           .rxpolarity11
		input  wire        rxpolarity12,              //           .rxpolarity12
		input  wire        rxpolarity13,              //           .rxpolarity13
		input  wire        rxpolarity14,              //           .rxpolarity14
		input  wire        rxpolarity15,              //           .rxpolarity15
		input  wire        txcompl8,                  //           .txcompl8
		input  wire        txcompl9,                  //           .txcompl9
		input  wire        txcompl10,                 //           .txcompl10
		input  wire        txcompl11,                 //           .txcompl11
		input  wire        txcompl12,                 //           .txcompl12
		input  wire        txcompl13,                 //           .txcompl13
		input  wire        txcompl14,                 //           .txcompl14
		input  wire        txcompl15,                 //           .txcompl15
		input  wire [31:0] txdata8,                   //           .txdata8
		input  wire [31:0] txdata9,                   //           .txdata9
		input  wire [31:0] txdata10,                  //           .txdata10
		input  wire [31:0] txdata11,                  //           .txdata11
		input  wire [31:0] txdata12,                  //           .txdata12
		input  wire [31:0] txdata13,                  //           .txdata13
		input  wire [31:0] txdata14,                  //           .txdata14
		input  wire [31:0] txdata15,                  //           .txdata15
		input  wire [3:0]  txdatak8,                  //           .txdatak8
		input  wire [3:0]  txdatak9,                  //           .txdatak9
		input  wire [3:0]  txdatak10,                 //           .txdatak10
		input  wire [3:0]  txdatak11,                 //           .txdatak11
		input  wire [3:0]  txdatak12,                 //           .txdatak12
		input  wire [3:0]  txdatak13,                 //           .txdatak13
		input  wire [3:0]  txdatak14,                 //           .txdatak14
		input  wire [3:0]  txdatak15,                 //           .txdatak15
		input  wire        txdetectrx8,               //           .txdetectrx8
		input  wire        txdetectrx9,               //           .txdetectrx9
		input  wire        txdetectrx10,              //           .txdetectrx10
		input  wire        txdetectrx11,              //           .txdetectrx11
		input  wire        txdetectrx12,              //           .txdetectrx12
		input  wire        txdetectrx13,              //           .txdetectrx13
		input  wire        txdetectrx14,              //           .txdetectrx14
		input  wire        txdetectrx15,              //           .txdetectrx15
		input  wire        txelecidle8,               //           .txelecidle8
		input  wire        txelecidle9,               //           .txelecidle9
		input  wire        txelecidle10,              //           .txelecidle10
		input  wire        txelecidle11,              //           .txelecidle11
		input  wire        txelecidle12,              //           .txelecidle12
		input  wire        txelecidle13,              //           .txelecidle13
		input  wire        txelecidle14,              //           .txelecidle14
		input  wire        txelecidle15,              //           .txelecidle15
		input  wire        txdeemph8,                 //           .txdeemph8
		input  wire        txdeemph9,                 //           .txdeemph9
		input  wire        txdeemph10,                //           .txdeemph10
		input  wire        txdeemph11,                //           .txdeemph11
		input  wire        txdeemph12,                //           .txdeemph12
		input  wire        txdeemph13,                //           .txdeemph13
		input  wire        txdeemph14,                //           .txdeemph14
		input  wire        txdeemph15,                //           .txdeemph15
		input  wire [2:0]  txmargin8,                 //           .txmargin8
		input  wire [2:0]  txmargin9,                 //           .txmargin9
		input  wire [2:0]  txmargin10,                //           .txmargin10
		input  wire [2:0]  txmargin11,                //           .txmargin11
		input  wire [2:0]  txmargin12,                //           .txmargin12
		input  wire [2:0]  txmargin13,                //           .txmargin13
		input  wire [2:0]  txmargin14,                //           .txmargin14
		input  wire [2:0]  txmargin15,                //           .txmargin15
		input  wire        txswing8,                  //           .txswing8
		input  wire        txswing9,                  //           .txswing9
		input  wire        txswing10,                 //           .txswing10
		input  wire        txswing11,                 //           .txswing11
		input  wire        txswing12,                 //           .txswing12
		input  wire        txswing13,                 //           .txswing13
		input  wire        txswing14,                 //           .txswing14
		input  wire        txswing15,                 //           .txswing15
		output wire        phystatus8,                //           .phystatus8
		output wire        phystatus9,                //           .phystatus9
		output wire        phystatus10,               //           .phystatus10
		output wire        phystatus11,               //           .phystatus11
		output wire        phystatus12,               //           .phystatus12
		output wire        phystatus13,               //           .phystatus13
		output wire        phystatus14,               //           .phystatus14
		output wire        phystatus15,               //           .phystatus15
		output wire [31:0] rxdata8,                   //           .rxdata8
		output wire [31:0] rxdata9,                   //           .rxdata9
		output wire [31:0] rxdata10,                  //           .rxdata10
		output wire [31:0] rxdata11,                  //           .rxdata11
		output wire [31:0] rxdata12,                  //           .rxdata12
		output wire [31:0] rxdata13,                  //           .rxdata13
		output wire [31:0] rxdata14,                  //           .rxdata14
		output wire [31:0] rxdata15,                  //           .rxdata15
		output wire [3:0]  rxdatak8,                  //           .rxdatak8
		output wire [3:0]  rxdatak9,                  //           .rxdatak9
		output wire [3:0]  rxdatak10,                 //           .rxdatak10
		output wire [3:0]  rxdatak11,                 //           .rxdatak11
		output wire [3:0]  rxdatak12,                 //           .rxdatak12
		output wire [3:0]  rxdatak13,                 //           .rxdatak13
		output wire [3:0]  rxdatak14,                 //           .rxdatak14
		output wire [3:0]  rxdatak15,                 //           .rxdatak15
		output wire        rxelecidle8,               //           .rxelecidle8
		output wire        rxelecidle9,               //           .rxelecidle9
		output wire        rxelecidle10,              //           .rxelecidle10
		output wire        rxelecidle11,              //           .rxelecidle11
		output wire        rxelecidle12,              //           .rxelecidle12
		output wire        rxelecidle13,              //           .rxelecidle13
		output wire        rxelecidle14,              //           .rxelecidle14
		output wire        rxelecidle15,              //           .rxelecidle15
		output wire [2:0]  rxstatus8,                 //           .rxstatus8
		output wire [2:0]  rxstatus9,                 //           .rxstatus9
		output wire [2:0]  rxstatus10,                //           .rxstatus10
		output wire [2:0]  rxstatus11,                //           .rxstatus11
		output wire [2:0]  rxstatus12,                //           .rxstatus12
		output wire [2:0]  rxstatus13,                //           .rxstatus13
		output wire [2:0]  rxstatus14,                //           .rxstatus14
		output wire [2:0]  rxstatus15,                //           .rxstatus15
		output wire        rxvalid8,                  //           .rxvalid8
		output wire        rxvalid9,                  //           .rxvalid9
		output wire        rxvalid10,                 //           .rxvalid10
		output wire        rxvalid11,                 //           .rxvalid11
		output wire        rxvalid12,                 //           .rxvalid12
		output wire        rxvalid13,                 //           .rxvalid13
		output wire        rxvalid14,                 //           .rxvalid14
		output wire        rxvalid15,                 //           .rxvalid15
		output wire        rxdataskip8,               //           .rxdataskip8
		output wire        rxdataskip9,               //           .rxdataskip9
		output wire        rxdataskip10,              //           .rxdataskip10
		output wire        rxdataskip11,              //           .rxdataskip11
		output wire        rxdataskip12,              //           .rxdataskip12
		output wire        rxdataskip13,              //           .rxdataskip13
		output wire        rxdataskip14,              //           .rxdataskip14
		output wire        rxdataskip15,              //           .rxdataskip15
		output wire        rxblkst8,                  //           .rxblkst8
		output wire        rxblkst9,                  //           .rxblkst9
		output wire        rxblkst10,                 //           .rxblkst10
		output wire        rxblkst11,                 //           .rxblkst11
		output wire        rxblkst12,                 //           .rxblkst12
		output wire        rxblkst13,                 //           .rxblkst13
		output wire        rxblkst14,                 //           .rxblkst14
		output wire        rxblkst15,                 //           .rxblkst15
		output wire [1:0]  rxsynchd8,                 //           .rxsynchd8
		output wire [1:0]  rxsynchd9,                 //           .rxsynchd9
		output wire [1:0]  rxsynchd10,                //           .rxsynchd10
		output wire [1:0]  rxsynchd11,                //           .rxsynchd11
		output wire [1:0]  rxsynchd12,                //           .rxsynchd12
		output wire [1:0]  rxsynchd13,                //           .rxsynchd13
		output wire [1:0]  rxsynchd14,                //           .rxsynchd14
		output wire [1:0]  rxsynchd15,                //           .rxsynchd15
		input  wire [17:0] currentcoeff8,             //           .currentcoeff8
		input  wire [17:0] currentcoeff9,             //           .currentcoeff9
		input  wire [17:0] currentcoeff10,            //           .currentcoeff10
		input  wire [17:0] currentcoeff11,            //           .currentcoeff11
		input  wire [17:0] currentcoeff12,            //           .currentcoeff12
		input  wire [17:0] currentcoeff13,            //           .currentcoeff13
		input  wire [17:0] currentcoeff14,            //           .currentcoeff14
		input  wire [17:0] currentcoeff15,            //           .currentcoeff15
		input  wire [2:0]  currentrxpreset8,          //           .currentrxpreset8
		input  wire [2:0]  currentrxpreset9,          //           .currentrxpreset9
		input  wire [2:0]  currentrxpreset10,         //           .currentrxpreset10
		input  wire [2:0]  currentrxpreset11,         //           .currentrxpreset11
		input  wire [2:0]  currentrxpreset12,         //           .currentrxpreset12
		input  wire [2:0]  currentrxpreset13,         //           .currentrxpreset13
		input  wire [2:0]  currentrxpreset14,         //           .currentrxpreset14
		input  wire [2:0]  currentrxpreset15,         //           .currentrxpreset15
		input  wire [1:0]  txsynchd8,                 //           .txsynchd8
		input  wire [1:0]  txsynchd9,                 //           .txsynchd9
		input  wire [1:0]  txsynchd10,                //           .txsynchd10
		input  wire [1:0]  txsynchd11,                //           .txsynchd11
		input  wire [1:0]  txsynchd12,                //           .txsynchd12
		input  wire [1:0]  txsynchd13,                //           .txsynchd13
		input  wire [1:0]  txsynchd14,                //           .txsynchd14
		input  wire [1:0]  txsynchd15,                //           .txsynchd15
		input  wire        txblkst8,                  //           .txblkst8
		input  wire        txblkst9,                  //           .txblkst9
		input  wire        txblkst10,                 //           .txblkst10
		input  wire        txblkst11,                 //           .txblkst11
		input  wire        txblkst12,                 //           .txblkst12
		input  wire        txblkst13,                 //           .txblkst13
		input  wire        txblkst14,                 //           .txblkst14
		input  wire        txblkst15,                 //           .txblkst15
		input  wire        txdataskip8,               //           .txdataskip8
		input  wire        txdataskip9,               //           .txdataskip9
		input  wire        txdataskip10,              //           .txdataskip10
		input  wire        txdataskip11,              //           .txdataskip11
		input  wire        txdataskip12,              //           .txdataskip12
		input  wire        txdataskip13,              //           .txdataskip13
		input  wire        txdataskip14,              //           .txdataskip14
		input  wire        txdataskip15,              //           .txdataskip15
		input  wire [1:0]  rate8,                     //           .rate8
		input  wire [1:0]  rate9,                     //           .rate9
		input  wire [1:0]  rate10,                    //           .rate10
		input  wire [1:0]  rate11,                    //           .rate11
		input  wire [1:0]  rate12,                    //           .rate12
		input  wire [1:0]  rate13,                    //           .rate13
		input  wire [1:0]  rate14,                    //           .rate14
		input  wire [1:0]  rate15,                    //           .rate15
		output wire [66:0] test_in,                   //   hip_ctrl.test_in
		output wire        simu_mode_pipe,            //           .simu_mode_pipe
		output wire        npor,                      //       npor.npor
		output wire        pin_perst                  //           .pin_perst
	);

	altpcie_s10_tbed_hwtcl #(
		.lane_mask_hwtcl                      (lane_mask_hwtcl),
		.gen123_lane_rate_mode_hwtcl          ("Gen3 (8.0 Gbps)"),
		.port_type_hwtcl                      ("Root Port"),
		.pll_refclk_freq_hwtcl                (pll_refclk_freq_hwtcl),
		.apps_type_hwtcl                      (13),
		.serial_sim_hwtcl                     (serial_sim_hwtcl),
		.deemphasis_enable_hwtcl              (deemphasis_enable_hwtcl),
		.pld_clk_MHz                          (pld_clk_MHz),
		.millisecond_cycle_count_hwtcl        (millisecond_cycle_count_hwtcl),
		.use_crc_forwarding_hwtcl             (use_crc_forwarding_hwtcl),
		.ecrc_check_capable_hwtcl             (ecrc_check_capable_hwtcl),
		.ecrc_gen_capable_hwtcl               (ecrc_gen_capable_hwtcl),
		.bfm_drive_interface_clk_hwtcl        (bfm_drive_interface_clk_hwtcl),
		.bfm_drive_interface_npor_hwtcl       (bfm_drive_interface_npor_hwtcl),
		.bfm_drive_interface_pipe_hwtcl       (bfm_drive_interface_pipe_hwtcl),
		.bfm_drive_interface_control_hwtcl    (bfm_drive_interface_control_hwtcl),
		.select_example_design_sim_BFM_hwtcl  (select_example_design_sim_BFM_hwtcl),
		.enable_pipe32_phyip_ser_driver_hwtcl (enable_pipe32_phyip_ser_driver_hwtcl)
	) dut_pcie_tb (
		.rx_in0                    (rx_in0),                    //  output,   width = 1, hip_serial.rx_in0
		.rx_in1                    (rx_in1),                    //  output,   width = 1,           .rx_in1
		.rx_in2                    (rx_in2),                    //  output,   width = 1,           .rx_in2
		.rx_in3                    (rx_in3),                    //  output,   width = 1,           .rx_in3
		.rx_in4                    (rx_in4),                    //  output,   width = 1,           .rx_in4
		.rx_in5                    (rx_in5),                    //  output,   width = 1,           .rx_in5
		.rx_in6                    (rx_in6),                    //  output,   width = 1,           .rx_in6
		.rx_in7                    (rx_in7),                    //  output,   width = 1,           .rx_in7
		.rx_in8                    (rx_in8),                    //  output,   width = 1,           .rx_in8
		.rx_in9                    (rx_in9),                    //  output,   width = 1,           .rx_in9
		.rx_in10                   (rx_in10),                   //  output,   width = 1,           .rx_in10
		.rx_in11                   (rx_in11),                   //  output,   width = 1,           .rx_in11
		.rx_in12                   (rx_in12),                   //  output,   width = 1,           .rx_in12
		.rx_in13                   (rx_in13),                   //  output,   width = 1,           .rx_in13
		.rx_in14                   (rx_in14),                   //  output,   width = 1,           .rx_in14
		.rx_in15                   (rx_in15),                   //  output,   width = 1,           .rx_in15
		.tx_out0                   (tx_out0),                   //   input,   width = 1,           .tx_out0
		.tx_out1                   (tx_out1),                   //   input,   width = 1,           .tx_out1
		.tx_out2                   (tx_out2),                   //   input,   width = 1,           .tx_out2
		.tx_out3                   (tx_out3),                   //   input,   width = 1,           .tx_out3
		.tx_out4                   (tx_out4),                   //   input,   width = 1,           .tx_out4
		.tx_out5                   (tx_out5),                   //   input,   width = 1,           .tx_out5
		.tx_out6                   (tx_out6),                   //   input,   width = 1,           .tx_out6
		.tx_out7                   (tx_out7),                   //   input,   width = 1,           .tx_out7
		.tx_out8                   (tx_out8),                   //   input,   width = 1,           .tx_out8
		.tx_out9                   (tx_out9),                   //   input,   width = 1,           .tx_out9
		.tx_out10                  (tx_out10),                  //   input,   width = 1,           .tx_out10
		.tx_out11                  (tx_out11),                  //   input,   width = 1,           .tx_out11
		.tx_out12                  (tx_out12),                  //   input,   width = 1,           .tx_out12
		.tx_out13                  (tx_out13),                  //   input,   width = 1,           .tx_out13
		.tx_out14                  (tx_out14),                  //   input,   width = 1,           .tx_out14
		.tx_out15                  (tx_out15),                  //   input,   width = 1,           .tx_out15
		.refclk                    (refclk),                    //  output,   width = 1,     refclk.clk
		.sim_pipe_pclk_in          (sim_pipe_pclk_in),          //  output,   width = 1,   hip_pipe.sim_pipe_pclk_in
		.sim_pipe_mask_tx_pll_lock (sim_pipe_mask_tx_pll_lock), //  output,   width = 1,           .sim_pipe_mask_tx_pll_lock
		.sim_pipe_rate             (sim_pipe_rate),             //   input,   width = 2,           .sim_pipe_rate
		.sim_ltssmstate            (sim_ltssmstate),            //   input,   width = 6,           .sim_ltssmstate
		.dirfeedback0              (dirfeedback0),              //  output,   width = 6,           .dirfeedback0
		.dirfeedback1              (dirfeedback1),              //  output,   width = 6,           .dirfeedback1
		.dirfeedback2              (dirfeedback2),              //  output,   width = 6,           .dirfeedback2
		.dirfeedback3              (dirfeedback3),              //  output,   width = 6,           .dirfeedback3
		.dirfeedback4              (dirfeedback4),              //  output,   width = 6,           .dirfeedback4
		.dirfeedback5              (dirfeedback5),              //  output,   width = 6,           .dirfeedback5
		.dirfeedback6              (dirfeedback6),              //  output,   width = 6,           .dirfeedback6
		.dirfeedback7              (dirfeedback7),              //  output,   width = 6,           .dirfeedback7
		.rxeqeval0                 (rxeqeval0),                 //   input,   width = 1,           .rxeqeval0
		.rxeqeval1                 (rxeqeval1),                 //   input,   width = 1,           .rxeqeval1
		.rxeqeval2                 (rxeqeval2),                 //   input,   width = 1,           .rxeqeval2
		.rxeqeval3                 (rxeqeval3),                 //   input,   width = 1,           .rxeqeval3
		.rxeqeval4                 (rxeqeval4),                 //   input,   width = 1,           .rxeqeval4
		.rxeqeval5                 (rxeqeval5),                 //   input,   width = 1,           .rxeqeval5
		.rxeqeval6                 (rxeqeval6),                 //   input,   width = 1,           .rxeqeval6
		.rxeqeval7                 (rxeqeval7),                 //   input,   width = 1,           .rxeqeval7
		.rxeqinprogress0           (rxeqinprogress0),           //   input,   width = 1,           .rxeqinprogress0
		.rxeqinprogress1           (rxeqinprogress1),           //   input,   width = 1,           .rxeqinprogress1
		.rxeqinprogress2           (rxeqinprogress2),           //   input,   width = 1,           .rxeqinprogress2
		.rxeqinprogress3           (rxeqinprogress3),           //   input,   width = 1,           .rxeqinprogress3
		.rxeqinprogress4           (rxeqinprogress4),           //   input,   width = 1,           .rxeqinprogress4
		.rxeqinprogress5           (rxeqinprogress5),           //   input,   width = 1,           .rxeqinprogress5
		.rxeqinprogress6           (rxeqinprogress6),           //   input,   width = 1,           .rxeqinprogress6
		.rxeqinprogress7           (rxeqinprogress7),           //   input,   width = 1,           .rxeqinprogress7
		.invalidreq0               (invalidreq0),               //   input,   width = 1,           .invalidreq0
		.invalidreq1               (invalidreq1),               //   input,   width = 1,           .invalidreq1
		.invalidreq2               (invalidreq2),               //   input,   width = 1,           .invalidreq2
		.invalidreq3               (invalidreq3),               //   input,   width = 1,           .invalidreq3
		.invalidreq4               (invalidreq4),               //   input,   width = 1,           .invalidreq4
		.invalidreq5               (invalidreq5),               //   input,   width = 1,           .invalidreq5
		.invalidreq6               (invalidreq6),               //   input,   width = 1,           .invalidreq6
		.invalidreq7               (invalidreq7),               //   input,   width = 1,           .invalidreq7
		.powerdown0                (powerdown0),                //   input,   width = 2,           .powerdown0
		.powerdown1                (powerdown1),                //   input,   width = 2,           .powerdown1
		.powerdown2                (powerdown2),                //   input,   width = 2,           .powerdown2
		.powerdown3                (powerdown3),                //   input,   width = 2,           .powerdown3
		.powerdown4                (powerdown4),                //   input,   width = 2,           .powerdown4
		.powerdown5                (powerdown5),                //   input,   width = 2,           .powerdown5
		.powerdown6                (powerdown6),                //   input,   width = 2,           .powerdown6
		.powerdown7                (powerdown7),                //   input,   width = 2,           .powerdown7
		.rxpolarity0               (rxpolarity0),               //   input,   width = 1,           .rxpolarity0
		.rxpolarity1               (rxpolarity1),               //   input,   width = 1,           .rxpolarity1
		.rxpolarity2               (rxpolarity2),               //   input,   width = 1,           .rxpolarity2
		.rxpolarity3               (rxpolarity3),               //   input,   width = 1,           .rxpolarity3
		.rxpolarity4               (rxpolarity4),               //   input,   width = 1,           .rxpolarity4
		.rxpolarity5               (rxpolarity5),               //   input,   width = 1,           .rxpolarity5
		.rxpolarity6               (rxpolarity6),               //   input,   width = 1,           .rxpolarity6
		.rxpolarity7               (rxpolarity7),               //   input,   width = 1,           .rxpolarity7
		.txcompl0                  (txcompl0),                  //   input,   width = 1,           .txcompl0
		.txcompl1                  (txcompl1),                  //   input,   width = 1,           .txcompl1
		.txcompl2                  (txcompl2),                  //   input,   width = 1,           .txcompl2
		.txcompl3                  (txcompl3),                  //   input,   width = 1,           .txcompl3
		.txcompl4                  (txcompl4),                  //   input,   width = 1,           .txcompl4
		.txcompl5                  (txcompl5),                  //   input,   width = 1,           .txcompl5
		.txcompl6                  (txcompl6),                  //   input,   width = 1,           .txcompl6
		.txcompl7                  (txcompl7),                  //   input,   width = 1,           .txcompl7
		.txdata0                   (txdata0),                   //   input,  width = 32,           .txdata0
		.txdata1                   (txdata1),                   //   input,  width = 32,           .txdata1
		.txdata2                   (txdata2),                   //   input,  width = 32,           .txdata2
		.txdata3                   (txdata3),                   //   input,  width = 32,           .txdata3
		.txdata4                   (txdata4),                   //   input,  width = 32,           .txdata4
		.txdata5                   (txdata5),                   //   input,  width = 32,           .txdata5
		.txdata6                   (txdata6),                   //   input,  width = 32,           .txdata6
		.txdata7                   (txdata7),                   //   input,  width = 32,           .txdata7
		.txdatak0                  (txdatak0),                  //   input,   width = 4,           .txdatak0
		.txdatak1                  (txdatak1),                  //   input,   width = 4,           .txdatak1
		.txdatak2                  (txdatak2),                  //   input,   width = 4,           .txdatak2
		.txdatak3                  (txdatak3),                  //   input,   width = 4,           .txdatak3
		.txdatak4                  (txdatak4),                  //   input,   width = 4,           .txdatak4
		.txdatak5                  (txdatak5),                  //   input,   width = 4,           .txdatak5
		.txdatak6                  (txdatak6),                  //   input,   width = 4,           .txdatak6
		.txdatak7                  (txdatak7),                  //   input,   width = 4,           .txdatak7
		.txdetectrx0               (txdetectrx0),               //   input,   width = 1,           .txdetectrx0
		.txdetectrx1               (txdetectrx1),               //   input,   width = 1,           .txdetectrx1
		.txdetectrx2               (txdetectrx2),               //   input,   width = 1,           .txdetectrx2
		.txdetectrx3               (txdetectrx3),               //   input,   width = 1,           .txdetectrx3
		.txdetectrx4               (txdetectrx4),               //   input,   width = 1,           .txdetectrx4
		.txdetectrx5               (txdetectrx5),               //   input,   width = 1,           .txdetectrx5
		.txdetectrx6               (txdetectrx6),               //   input,   width = 1,           .txdetectrx6
		.txdetectrx7               (txdetectrx7),               //   input,   width = 1,           .txdetectrx7
		.txelecidle0               (txelecidle0),               //   input,   width = 1,           .txelecidle0
		.txelecidle1               (txelecidle1),               //   input,   width = 1,           .txelecidle1
		.txelecidle2               (txelecidle2),               //   input,   width = 1,           .txelecidle2
		.txelecidle3               (txelecidle3),               //   input,   width = 1,           .txelecidle3
		.txelecidle4               (txelecidle4),               //   input,   width = 1,           .txelecidle4
		.txelecidle5               (txelecidle5),               //   input,   width = 1,           .txelecidle5
		.txelecidle6               (txelecidle6),               //   input,   width = 1,           .txelecidle6
		.txelecidle7               (txelecidle7),               //   input,   width = 1,           .txelecidle7
		.txdeemph0                 (txdeemph0),                 //   input,   width = 1,           .txdeemph0
		.txdeemph1                 (txdeemph1),                 //   input,   width = 1,           .txdeemph1
		.txdeemph2                 (txdeemph2),                 //   input,   width = 1,           .txdeemph2
		.txdeemph3                 (txdeemph3),                 //   input,   width = 1,           .txdeemph3
		.txdeemph4                 (txdeemph4),                 //   input,   width = 1,           .txdeemph4
		.txdeemph5                 (txdeemph5),                 //   input,   width = 1,           .txdeemph5
		.txdeemph6                 (txdeemph6),                 //   input,   width = 1,           .txdeemph6
		.txdeemph7                 (txdeemph7),                 //   input,   width = 1,           .txdeemph7
		.txmargin0                 (txmargin0),                 //   input,   width = 3,           .txmargin0
		.txmargin1                 (txmargin1),                 //   input,   width = 3,           .txmargin1
		.txmargin2                 (txmargin2),                 //   input,   width = 3,           .txmargin2
		.txmargin3                 (txmargin3),                 //   input,   width = 3,           .txmargin3
		.txmargin4                 (txmargin4),                 //   input,   width = 3,           .txmargin4
		.txmargin5                 (txmargin5),                 //   input,   width = 3,           .txmargin5
		.txmargin6                 (txmargin6),                 //   input,   width = 3,           .txmargin6
		.txmargin7                 (txmargin7),                 //   input,   width = 3,           .txmargin7
		.txswing0                  (txswing0),                  //   input,   width = 1,           .txswing0
		.txswing1                  (txswing1),                  //   input,   width = 1,           .txswing1
		.txswing2                  (txswing2),                  //   input,   width = 1,           .txswing2
		.txswing3                  (txswing3),                  //   input,   width = 1,           .txswing3
		.txswing4                  (txswing4),                  //   input,   width = 1,           .txswing4
		.txswing5                  (txswing5),                  //   input,   width = 1,           .txswing5
		.txswing6                  (txswing6),                  //   input,   width = 1,           .txswing6
		.txswing7                  (txswing7),                  //   input,   width = 1,           .txswing7
		.phystatus0                (phystatus0),                //  output,   width = 1,           .phystatus0
		.phystatus1                (phystatus1),                //  output,   width = 1,           .phystatus1
		.phystatus2                (phystatus2),                //  output,   width = 1,           .phystatus2
		.phystatus3                (phystatus3),                //  output,   width = 1,           .phystatus3
		.phystatus4                (phystatus4),                //  output,   width = 1,           .phystatus4
		.phystatus5                (phystatus5),                //  output,   width = 1,           .phystatus5
		.phystatus6                (phystatus6),                //  output,   width = 1,           .phystatus6
		.phystatus7                (phystatus7),                //  output,   width = 1,           .phystatus7
		.rxdata0                   (rxdata0),                   //  output,  width = 32,           .rxdata0
		.rxdata1                   (rxdata1),                   //  output,  width = 32,           .rxdata1
		.rxdata2                   (rxdata2),                   //  output,  width = 32,           .rxdata2
		.rxdata3                   (rxdata3),                   //  output,  width = 32,           .rxdata3
		.rxdata4                   (rxdata4),                   //  output,  width = 32,           .rxdata4
		.rxdata5                   (rxdata5),                   //  output,  width = 32,           .rxdata5
		.rxdata6                   (rxdata6),                   //  output,  width = 32,           .rxdata6
		.rxdata7                   (rxdata7),                   //  output,  width = 32,           .rxdata7
		.rxdatak0                  (rxdatak0),                  //  output,   width = 4,           .rxdatak0
		.rxdatak1                  (rxdatak1),                  //  output,   width = 4,           .rxdatak1
		.rxdatak2                  (rxdatak2),                  //  output,   width = 4,           .rxdatak2
		.rxdatak3                  (rxdatak3),                  //  output,   width = 4,           .rxdatak3
		.rxdatak4                  (rxdatak4),                  //  output,   width = 4,           .rxdatak4
		.rxdatak5                  (rxdatak5),                  //  output,   width = 4,           .rxdatak5
		.rxdatak6                  (rxdatak6),                  //  output,   width = 4,           .rxdatak6
		.rxdatak7                  (rxdatak7),                  //  output,   width = 4,           .rxdatak7
		.rxelecidle0               (rxelecidle0),               //  output,   width = 1,           .rxelecidle0
		.rxelecidle1               (rxelecidle1),               //  output,   width = 1,           .rxelecidle1
		.rxelecidle2               (rxelecidle2),               //  output,   width = 1,           .rxelecidle2
		.rxelecidle3               (rxelecidle3),               //  output,   width = 1,           .rxelecidle3
		.rxelecidle4               (rxelecidle4),               //  output,   width = 1,           .rxelecidle4
		.rxelecidle5               (rxelecidle5),               //  output,   width = 1,           .rxelecidle5
		.rxelecidle6               (rxelecidle6),               //  output,   width = 1,           .rxelecidle6
		.rxelecidle7               (rxelecidle7),               //  output,   width = 1,           .rxelecidle7
		.rxstatus0                 (rxstatus0),                 //  output,   width = 3,           .rxstatus0
		.rxstatus1                 (rxstatus1),                 //  output,   width = 3,           .rxstatus1
		.rxstatus2                 (rxstatus2),                 //  output,   width = 3,           .rxstatus2
		.rxstatus3                 (rxstatus3),                 //  output,   width = 3,           .rxstatus3
		.rxstatus4                 (rxstatus4),                 //  output,   width = 3,           .rxstatus4
		.rxstatus5                 (rxstatus5),                 //  output,   width = 3,           .rxstatus5
		.rxstatus6                 (rxstatus6),                 //  output,   width = 3,           .rxstatus6
		.rxstatus7                 (rxstatus7),                 //  output,   width = 3,           .rxstatus7
		.rxvalid0                  (rxvalid0),                  //  output,   width = 1,           .rxvalid0
		.rxvalid1                  (rxvalid1),                  //  output,   width = 1,           .rxvalid1
		.rxvalid2                  (rxvalid2),                  //  output,   width = 1,           .rxvalid2
		.rxvalid3                  (rxvalid3),                  //  output,   width = 1,           .rxvalid3
		.rxvalid4                  (rxvalid4),                  //  output,   width = 1,           .rxvalid4
		.rxvalid5                  (rxvalid5),                  //  output,   width = 1,           .rxvalid5
		.rxvalid6                  (rxvalid6),                  //  output,   width = 1,           .rxvalid6
		.rxvalid7                  (rxvalid7),                  //  output,   width = 1,           .rxvalid7
		.rxdataskip0               (rxdataskip0),               //  output,   width = 1,           .rxdataskip0
		.rxdataskip1               (rxdataskip1),               //  output,   width = 1,           .rxdataskip1
		.rxdataskip2               (rxdataskip2),               //  output,   width = 1,           .rxdataskip2
		.rxdataskip3               (rxdataskip3),               //  output,   width = 1,           .rxdataskip3
		.rxdataskip4               (rxdataskip4),               //  output,   width = 1,           .rxdataskip4
		.rxdataskip5               (rxdataskip5),               //  output,   width = 1,           .rxdataskip5
		.rxdataskip6               (rxdataskip6),               //  output,   width = 1,           .rxdataskip6
		.rxdataskip7               (rxdataskip7),               //  output,   width = 1,           .rxdataskip7
		.rxblkst0                  (rxblkst0),                  //  output,   width = 1,           .rxblkst0
		.rxblkst1                  (rxblkst1),                  //  output,   width = 1,           .rxblkst1
		.rxblkst2                  (rxblkst2),                  //  output,   width = 1,           .rxblkst2
		.rxblkst3                  (rxblkst3),                  //  output,   width = 1,           .rxblkst3
		.rxblkst4                  (rxblkst4),                  //  output,   width = 1,           .rxblkst4
		.rxblkst5                  (rxblkst5),                  //  output,   width = 1,           .rxblkst5
		.rxblkst6                  (rxblkst6),                  //  output,   width = 1,           .rxblkst6
		.rxblkst7                  (rxblkst7),                  //  output,   width = 1,           .rxblkst7
		.rxsynchd0                 (rxsynchd0),                 //  output,   width = 2,           .rxsynchd0
		.rxsynchd1                 (rxsynchd1),                 //  output,   width = 2,           .rxsynchd1
		.rxsynchd2                 (rxsynchd2),                 //  output,   width = 2,           .rxsynchd2
		.rxsynchd3                 (rxsynchd3),                 //  output,   width = 2,           .rxsynchd3
		.rxsynchd4                 (rxsynchd4),                 //  output,   width = 2,           .rxsynchd4
		.rxsynchd5                 (rxsynchd5),                 //  output,   width = 2,           .rxsynchd5
		.rxsynchd6                 (rxsynchd6),                 //  output,   width = 2,           .rxsynchd6
		.rxsynchd7                 (rxsynchd7),                 //  output,   width = 2,           .rxsynchd7
		.currentcoeff0             (currentcoeff0),             //   input,  width = 18,           .currentcoeff0
		.currentcoeff1             (currentcoeff1),             //   input,  width = 18,           .currentcoeff1
		.currentcoeff2             (currentcoeff2),             //   input,  width = 18,           .currentcoeff2
		.currentcoeff3             (currentcoeff3),             //   input,  width = 18,           .currentcoeff3
		.currentcoeff4             (currentcoeff4),             //   input,  width = 18,           .currentcoeff4
		.currentcoeff5             (currentcoeff5),             //   input,  width = 18,           .currentcoeff5
		.currentcoeff6             (currentcoeff6),             //   input,  width = 18,           .currentcoeff6
		.currentcoeff7             (currentcoeff7),             //   input,  width = 18,           .currentcoeff7
		.currentrxpreset0          (currentrxpreset0),          //   input,   width = 3,           .currentrxpreset0
		.currentrxpreset1          (currentrxpreset1),          //   input,   width = 3,           .currentrxpreset1
		.currentrxpreset2          (currentrxpreset2),          //   input,   width = 3,           .currentrxpreset2
		.currentrxpreset3          (currentrxpreset3),          //   input,   width = 3,           .currentrxpreset3
		.currentrxpreset4          (currentrxpreset4),          //   input,   width = 3,           .currentrxpreset4
		.currentrxpreset5          (currentrxpreset5),          //   input,   width = 3,           .currentrxpreset5
		.currentrxpreset6          (currentrxpreset6),          //   input,   width = 3,           .currentrxpreset6
		.currentrxpreset7          (currentrxpreset7),          //   input,   width = 3,           .currentrxpreset7
		.txsynchd0                 (txsynchd0),                 //   input,   width = 2,           .txsynchd0
		.txsynchd1                 (txsynchd1),                 //   input,   width = 2,           .txsynchd1
		.txsynchd2                 (txsynchd2),                 //   input,   width = 2,           .txsynchd2
		.txsynchd3                 (txsynchd3),                 //   input,   width = 2,           .txsynchd3
		.txsynchd4                 (txsynchd4),                 //   input,   width = 2,           .txsynchd4
		.txsynchd5                 (txsynchd5),                 //   input,   width = 2,           .txsynchd5
		.txsynchd6                 (txsynchd6),                 //   input,   width = 2,           .txsynchd6
		.txsynchd7                 (txsynchd7),                 //   input,   width = 2,           .txsynchd7
		.txblkst0                  (txblkst0),                  //   input,   width = 1,           .txblkst0
		.txblkst1                  (txblkst1),                  //   input,   width = 1,           .txblkst1
		.txblkst2                  (txblkst2),                  //   input,   width = 1,           .txblkst2
		.txblkst3                  (txblkst3),                  //   input,   width = 1,           .txblkst3
		.txblkst4                  (txblkst4),                  //   input,   width = 1,           .txblkst4
		.txblkst5                  (txblkst5),                  //   input,   width = 1,           .txblkst5
		.txblkst6                  (txblkst6),                  //   input,   width = 1,           .txblkst6
		.txblkst7                  (txblkst7),                  //   input,   width = 1,           .txblkst7
		.txdataskip0               (txdataskip0),               //   input,   width = 1,           .txdataskip0
		.txdataskip1               (txdataskip1),               //   input,   width = 1,           .txdataskip1
		.txdataskip2               (txdataskip2),               //   input,   width = 1,           .txdataskip2
		.txdataskip3               (txdataskip3),               //   input,   width = 1,           .txdataskip3
		.txdataskip4               (txdataskip4),               //   input,   width = 1,           .txdataskip4
		.txdataskip5               (txdataskip5),               //   input,   width = 1,           .txdataskip5
		.txdataskip6               (txdataskip6),               //   input,   width = 1,           .txdataskip6
		.txdataskip7               (txdataskip7),               //   input,   width = 1,           .txdataskip7
		.rate0                     (rate0),                     //   input,   width = 2,           .rate0
		.rate1                     (rate1),                     //   input,   width = 2,           .rate1
		.rate2                     (rate2),                     //   input,   width = 2,           .rate2
		.rate3                     (rate3),                     //   input,   width = 2,           .rate3
		.rate4                     (rate4),                     //   input,   width = 2,           .rate4
		.rate5                     (rate5),                     //   input,   width = 2,           .rate5
		.rate6                     (rate6),                     //   input,   width = 2,           .rate6
		.rate7                     (rate7),                     //   input,   width = 2,           .rate7
		.dirfeedback8              (dirfeedback8),              //  output,   width = 6,           .dirfeedback8
		.dirfeedback9              (dirfeedback9),              //  output,   width = 6,           .dirfeedback9
		.dirfeedback10             (dirfeedback10),             //  output,   width = 6,           .dirfeedback10
		.dirfeedback11             (dirfeedback11),             //  output,   width = 6,           .dirfeedback11
		.dirfeedback12             (dirfeedback12),             //  output,   width = 6,           .dirfeedback12
		.dirfeedback13             (dirfeedback13),             //  output,   width = 6,           .dirfeedback13
		.dirfeedback14             (dirfeedback14),             //  output,   width = 6,           .dirfeedback14
		.dirfeedback15             (dirfeedback15),             //  output,   width = 6,           .dirfeedback15
		.rxeqeval8                 (rxeqeval8),                 //   input,   width = 1,           .rxeqeval8
		.rxeqeval9                 (rxeqeval9),                 //   input,   width = 1,           .rxeqeval9
		.rxeqeval10                (rxeqeval10),                //   input,   width = 1,           .rxeqeval10
		.rxeqeval11                (rxeqeval11),                //   input,   width = 1,           .rxeqeval11
		.rxeqeval12                (rxeqeval12),                //   input,   width = 1,           .rxeqeval12
		.rxeqeval13                (rxeqeval13),                //   input,   width = 1,           .rxeqeval13
		.rxeqeval14                (rxeqeval14),                //   input,   width = 1,           .rxeqeval14
		.rxeqeval15                (rxeqeval15),                //   input,   width = 1,           .rxeqeval15
		.rxeqinprogress8           (rxeqinprogress8),           //   input,   width = 1,           .rxeqinprogress8
		.rxeqinprogress9           (rxeqinprogress9),           //   input,   width = 1,           .rxeqinprogress9
		.rxeqinprogress10          (rxeqinprogress10),          //   input,   width = 1,           .rxeqinprogress10
		.rxeqinprogress11          (rxeqinprogress11),          //   input,   width = 1,           .rxeqinprogress11
		.rxeqinprogress12          (rxeqinprogress12),          //   input,   width = 1,           .rxeqinprogress12
		.rxeqinprogress13          (rxeqinprogress13),          //   input,   width = 1,           .rxeqinprogress13
		.rxeqinprogress14          (rxeqinprogress14),          //   input,   width = 1,           .rxeqinprogress14
		.rxeqinprogress15          (rxeqinprogress15),          //   input,   width = 1,           .rxeqinprogress15
		.invalidreq8               (invalidreq8),               //   input,   width = 1,           .invalidreq8
		.invalidreq9               (invalidreq9),               //   input,   width = 1,           .invalidreq9
		.invalidreq10              (invalidreq10),              //   input,   width = 1,           .invalidreq10
		.invalidreq11              (invalidreq11),              //   input,   width = 1,           .invalidreq11
		.invalidreq12              (invalidreq12),              //   input,   width = 1,           .invalidreq12
		.invalidreq13              (invalidreq13),              //   input,   width = 1,           .invalidreq13
		.invalidreq14              (invalidreq14),              //   input,   width = 1,           .invalidreq14
		.invalidreq15              (invalidreq15),              //   input,   width = 1,           .invalidreq15
		.powerdown8                (powerdown8),                //   input,   width = 2,           .powerdown8
		.powerdown9                (powerdown9),                //   input,   width = 2,           .powerdown9
		.powerdown10               (powerdown10),               //   input,   width = 2,           .powerdown10
		.powerdown11               (powerdown11),               //   input,   width = 2,           .powerdown11
		.powerdown12               (powerdown12),               //   input,   width = 2,           .powerdown12
		.powerdown13               (powerdown13),               //   input,   width = 2,           .powerdown13
		.powerdown14               (powerdown14),               //   input,   width = 2,           .powerdown14
		.powerdown15               (powerdown15),               //   input,   width = 2,           .powerdown15
		.rxpolarity8               (rxpolarity8),               //   input,   width = 1,           .rxpolarity8
		.rxpolarity9               (rxpolarity9),               //   input,   width = 1,           .rxpolarity9
		.rxpolarity10              (rxpolarity10),              //   input,   width = 1,           .rxpolarity10
		.rxpolarity11              (rxpolarity11),              //   input,   width = 1,           .rxpolarity11
		.rxpolarity12              (rxpolarity12),              //   input,   width = 1,           .rxpolarity12
		.rxpolarity13              (rxpolarity13),              //   input,   width = 1,           .rxpolarity13
		.rxpolarity14              (rxpolarity14),              //   input,   width = 1,           .rxpolarity14
		.rxpolarity15              (rxpolarity15),              //   input,   width = 1,           .rxpolarity15
		.txcompl8                  (txcompl8),                  //   input,   width = 1,           .txcompl8
		.txcompl9                  (txcompl9),                  //   input,   width = 1,           .txcompl9
		.txcompl10                 (txcompl10),                 //   input,   width = 1,           .txcompl10
		.txcompl11                 (txcompl11),                 //   input,   width = 1,           .txcompl11
		.txcompl12                 (txcompl12),                 //   input,   width = 1,           .txcompl12
		.txcompl13                 (txcompl13),                 //   input,   width = 1,           .txcompl13
		.txcompl14                 (txcompl14),                 //   input,   width = 1,           .txcompl14
		.txcompl15                 (txcompl15),                 //   input,   width = 1,           .txcompl15
		.txdata8                   (txdata8),                   //   input,  width = 32,           .txdata8
		.txdata9                   (txdata9),                   //   input,  width = 32,           .txdata9
		.txdata10                  (txdata10),                  //   input,  width = 32,           .txdata10
		.txdata11                  (txdata11),                  //   input,  width = 32,           .txdata11
		.txdata12                  (txdata12),                  //   input,  width = 32,           .txdata12
		.txdata13                  (txdata13),                  //   input,  width = 32,           .txdata13
		.txdata14                  (txdata14),                  //   input,  width = 32,           .txdata14
		.txdata15                  (txdata15),                  //   input,  width = 32,           .txdata15
		.txdatak8                  (txdatak8),                  //   input,   width = 4,           .txdatak8
		.txdatak9                  (txdatak9),                  //   input,   width = 4,           .txdatak9
		.txdatak10                 (txdatak10),                 //   input,   width = 4,           .txdatak10
		.txdatak11                 (txdatak11),                 //   input,   width = 4,           .txdatak11
		.txdatak12                 (txdatak12),                 //   input,   width = 4,           .txdatak12
		.txdatak13                 (txdatak13),                 //   input,   width = 4,           .txdatak13
		.txdatak14                 (txdatak14),                 //   input,   width = 4,           .txdatak14
		.txdatak15                 (txdatak15),                 //   input,   width = 4,           .txdatak15
		.txdetectrx8               (txdetectrx8),               //   input,   width = 1,           .txdetectrx8
		.txdetectrx9               (txdetectrx9),               //   input,   width = 1,           .txdetectrx9
		.txdetectrx10              (txdetectrx10),              //   input,   width = 1,           .txdetectrx10
		.txdetectrx11              (txdetectrx11),              //   input,   width = 1,           .txdetectrx11
		.txdetectrx12              (txdetectrx12),              //   input,   width = 1,           .txdetectrx12
		.txdetectrx13              (txdetectrx13),              //   input,   width = 1,           .txdetectrx13
		.txdetectrx14              (txdetectrx14),              //   input,   width = 1,           .txdetectrx14
		.txdetectrx15              (txdetectrx15),              //   input,   width = 1,           .txdetectrx15
		.txelecidle8               (txelecidle8),               //   input,   width = 1,           .txelecidle8
		.txelecidle9               (txelecidle9),               //   input,   width = 1,           .txelecidle9
		.txelecidle10              (txelecidle10),              //   input,   width = 1,           .txelecidle10
		.txelecidle11              (txelecidle11),              //   input,   width = 1,           .txelecidle11
		.txelecidle12              (txelecidle12),              //   input,   width = 1,           .txelecidle12
		.txelecidle13              (txelecidle13),              //   input,   width = 1,           .txelecidle13
		.txelecidle14              (txelecidle14),              //   input,   width = 1,           .txelecidle14
		.txelecidle15              (txelecidle15),              //   input,   width = 1,           .txelecidle15
		.txdeemph8                 (txdeemph8),                 //   input,   width = 1,           .txdeemph8
		.txdeemph9                 (txdeemph9),                 //   input,   width = 1,           .txdeemph9
		.txdeemph10                (txdeemph10),                //   input,   width = 1,           .txdeemph10
		.txdeemph11                (txdeemph11),                //   input,   width = 1,           .txdeemph11
		.txdeemph12                (txdeemph12),                //   input,   width = 1,           .txdeemph12
		.txdeemph13                (txdeemph13),                //   input,   width = 1,           .txdeemph13
		.txdeemph14                (txdeemph14),                //   input,   width = 1,           .txdeemph14
		.txdeemph15                (txdeemph15),                //   input,   width = 1,           .txdeemph15
		.txmargin8                 (txmargin8),                 //   input,   width = 3,           .txmargin8
		.txmargin9                 (txmargin9),                 //   input,   width = 3,           .txmargin9
		.txmargin10                (txmargin10),                //   input,   width = 3,           .txmargin10
		.txmargin11                (txmargin11),                //   input,   width = 3,           .txmargin11
		.txmargin12                (txmargin12),                //   input,   width = 3,           .txmargin12
		.txmargin13                (txmargin13),                //   input,   width = 3,           .txmargin13
		.txmargin14                (txmargin14),                //   input,   width = 3,           .txmargin14
		.txmargin15                (txmargin15),                //   input,   width = 3,           .txmargin15
		.txswing8                  (txswing8),                  //   input,   width = 1,           .txswing8
		.txswing9                  (txswing9),                  //   input,   width = 1,           .txswing9
		.txswing10                 (txswing10),                 //   input,   width = 1,           .txswing10
		.txswing11                 (txswing11),                 //   input,   width = 1,           .txswing11
		.txswing12                 (txswing12),                 //   input,   width = 1,           .txswing12
		.txswing13                 (txswing13),                 //   input,   width = 1,           .txswing13
		.txswing14                 (txswing14),                 //   input,   width = 1,           .txswing14
		.txswing15                 (txswing15),                 //   input,   width = 1,           .txswing15
		.phystatus8                (phystatus8),                //  output,   width = 1,           .phystatus8
		.phystatus9                (phystatus9),                //  output,   width = 1,           .phystatus9
		.phystatus10               (phystatus10),               //  output,   width = 1,           .phystatus10
		.phystatus11               (phystatus11),               //  output,   width = 1,           .phystatus11
		.phystatus12               (phystatus12),               //  output,   width = 1,           .phystatus12
		.phystatus13               (phystatus13),               //  output,   width = 1,           .phystatus13
		.phystatus14               (phystatus14),               //  output,   width = 1,           .phystatus14
		.phystatus15               (phystatus15),               //  output,   width = 1,           .phystatus15
		.rxdata8                   (rxdata8),                   //  output,  width = 32,           .rxdata8
		.rxdata9                   (rxdata9),                   //  output,  width = 32,           .rxdata9
		.rxdata10                  (rxdata10),                  //  output,  width = 32,           .rxdata10
		.rxdata11                  (rxdata11),                  //  output,  width = 32,           .rxdata11
		.rxdata12                  (rxdata12),                  //  output,  width = 32,           .rxdata12
		.rxdata13                  (rxdata13),                  //  output,  width = 32,           .rxdata13
		.rxdata14                  (rxdata14),                  //  output,  width = 32,           .rxdata14
		.rxdata15                  (rxdata15),                  //  output,  width = 32,           .rxdata15
		.rxdatak8                  (rxdatak8),                  //  output,   width = 4,           .rxdatak8
		.rxdatak9                  (rxdatak9),                  //  output,   width = 4,           .rxdatak9
		.rxdatak10                 (rxdatak10),                 //  output,   width = 4,           .rxdatak10
		.rxdatak11                 (rxdatak11),                 //  output,   width = 4,           .rxdatak11
		.rxdatak12                 (rxdatak12),                 //  output,   width = 4,           .rxdatak12
		.rxdatak13                 (rxdatak13),                 //  output,   width = 4,           .rxdatak13
		.rxdatak14                 (rxdatak14),                 //  output,   width = 4,           .rxdatak14
		.rxdatak15                 (rxdatak15),                 //  output,   width = 4,           .rxdatak15
		.rxelecidle8               (rxelecidle8),               //  output,   width = 1,           .rxelecidle8
		.rxelecidle9               (rxelecidle9),               //  output,   width = 1,           .rxelecidle9
		.rxelecidle10              (rxelecidle10),              //  output,   width = 1,           .rxelecidle10
		.rxelecidle11              (rxelecidle11),              //  output,   width = 1,           .rxelecidle11
		.rxelecidle12              (rxelecidle12),              //  output,   width = 1,           .rxelecidle12
		.rxelecidle13              (rxelecidle13),              //  output,   width = 1,           .rxelecidle13
		.rxelecidle14              (rxelecidle14),              //  output,   width = 1,           .rxelecidle14
		.rxelecidle15              (rxelecidle15),              //  output,   width = 1,           .rxelecidle15
		.rxstatus8                 (rxstatus8),                 //  output,   width = 3,           .rxstatus8
		.rxstatus9                 (rxstatus9),                 //  output,   width = 3,           .rxstatus9
		.rxstatus10                (rxstatus10),                //  output,   width = 3,           .rxstatus10
		.rxstatus11                (rxstatus11),                //  output,   width = 3,           .rxstatus11
		.rxstatus12                (rxstatus12),                //  output,   width = 3,           .rxstatus12
		.rxstatus13                (rxstatus13),                //  output,   width = 3,           .rxstatus13
		.rxstatus14                (rxstatus14),                //  output,   width = 3,           .rxstatus14
		.rxstatus15                (rxstatus15),                //  output,   width = 3,           .rxstatus15
		.rxvalid8                  (rxvalid8),                  //  output,   width = 1,           .rxvalid8
		.rxvalid9                  (rxvalid9),                  //  output,   width = 1,           .rxvalid9
		.rxvalid10                 (rxvalid10),                 //  output,   width = 1,           .rxvalid10
		.rxvalid11                 (rxvalid11),                 //  output,   width = 1,           .rxvalid11
		.rxvalid12                 (rxvalid12),                 //  output,   width = 1,           .rxvalid12
		.rxvalid13                 (rxvalid13),                 //  output,   width = 1,           .rxvalid13
		.rxvalid14                 (rxvalid14),                 //  output,   width = 1,           .rxvalid14
		.rxvalid15                 (rxvalid15),                 //  output,   width = 1,           .rxvalid15
		.rxdataskip8               (rxdataskip8),               //  output,   width = 1,           .rxdataskip8
		.rxdataskip9               (rxdataskip9),               //  output,   width = 1,           .rxdataskip9
		.rxdataskip10              (rxdataskip10),              //  output,   width = 1,           .rxdataskip10
		.rxdataskip11              (rxdataskip11),              //  output,   width = 1,           .rxdataskip11
		.rxdataskip12              (rxdataskip12),              //  output,   width = 1,           .rxdataskip12
		.rxdataskip13              (rxdataskip13),              //  output,   width = 1,           .rxdataskip13
		.rxdataskip14              (rxdataskip14),              //  output,   width = 1,           .rxdataskip14
		.rxdataskip15              (rxdataskip15),              //  output,   width = 1,           .rxdataskip15
		.rxblkst8                  (rxblkst8),                  //  output,   width = 1,           .rxblkst8
		.rxblkst9                  (rxblkst9),                  //  output,   width = 1,           .rxblkst9
		.rxblkst10                 (rxblkst10),                 //  output,   width = 1,           .rxblkst10
		.rxblkst11                 (rxblkst11),                 //  output,   width = 1,           .rxblkst11
		.rxblkst12                 (rxblkst12),                 //  output,   width = 1,           .rxblkst12
		.rxblkst13                 (rxblkst13),                 //  output,   width = 1,           .rxblkst13
		.rxblkst14                 (rxblkst14),                 //  output,   width = 1,           .rxblkst14
		.rxblkst15                 (rxblkst15),                 //  output,   width = 1,           .rxblkst15
		.rxsynchd8                 (rxsynchd8),                 //  output,   width = 2,           .rxsynchd8
		.rxsynchd9                 (rxsynchd9),                 //  output,   width = 2,           .rxsynchd9
		.rxsynchd10                (rxsynchd10),                //  output,   width = 2,           .rxsynchd10
		.rxsynchd11                (rxsynchd11),                //  output,   width = 2,           .rxsynchd11
		.rxsynchd12                (rxsynchd12),                //  output,   width = 2,           .rxsynchd12
		.rxsynchd13                (rxsynchd13),                //  output,   width = 2,           .rxsynchd13
		.rxsynchd14                (rxsynchd14),                //  output,   width = 2,           .rxsynchd14
		.rxsynchd15                (rxsynchd15),                //  output,   width = 2,           .rxsynchd15
		.currentcoeff8             (currentcoeff8),             //   input,  width = 18,           .currentcoeff8
		.currentcoeff9             (currentcoeff9),             //   input,  width = 18,           .currentcoeff9
		.currentcoeff10            (currentcoeff10),            //   input,  width = 18,           .currentcoeff10
		.currentcoeff11            (currentcoeff11),            //   input,  width = 18,           .currentcoeff11
		.currentcoeff12            (currentcoeff12),            //   input,  width = 18,           .currentcoeff12
		.currentcoeff13            (currentcoeff13),            //   input,  width = 18,           .currentcoeff13
		.currentcoeff14            (currentcoeff14),            //   input,  width = 18,           .currentcoeff14
		.currentcoeff15            (currentcoeff15),            //   input,  width = 18,           .currentcoeff15
		.currentrxpreset8          (currentrxpreset8),          //   input,   width = 3,           .currentrxpreset8
		.currentrxpreset9          (currentrxpreset9),          //   input,   width = 3,           .currentrxpreset9
		.currentrxpreset10         (currentrxpreset10),         //   input,   width = 3,           .currentrxpreset10
		.currentrxpreset11         (currentrxpreset11),         //   input,   width = 3,           .currentrxpreset11
		.currentrxpreset12         (currentrxpreset12),         //   input,   width = 3,           .currentrxpreset12
		.currentrxpreset13         (currentrxpreset13),         //   input,   width = 3,           .currentrxpreset13
		.currentrxpreset14         (currentrxpreset14),         //   input,   width = 3,           .currentrxpreset14
		.currentrxpreset15         (currentrxpreset15),         //   input,   width = 3,           .currentrxpreset15
		.txsynchd8                 (txsynchd8),                 //   input,   width = 2,           .txsynchd8
		.txsynchd9                 (txsynchd9),                 //   input,   width = 2,           .txsynchd9
		.txsynchd10                (txsynchd10),                //   input,   width = 2,           .txsynchd10
		.txsynchd11                (txsynchd11),                //   input,   width = 2,           .txsynchd11
		.txsynchd12                (txsynchd12),                //   input,   width = 2,           .txsynchd12
		.txsynchd13                (txsynchd13),                //   input,   width = 2,           .txsynchd13
		.txsynchd14                (txsynchd14),                //   input,   width = 2,           .txsynchd14
		.txsynchd15                (txsynchd15),                //   input,   width = 2,           .txsynchd15
		.txblkst8                  (txblkst8),                  //   input,   width = 1,           .txblkst8
		.txblkst9                  (txblkst9),                  //   input,   width = 1,           .txblkst9
		.txblkst10                 (txblkst10),                 //   input,   width = 1,           .txblkst10
		.txblkst11                 (txblkst11),                 //   input,   width = 1,           .txblkst11
		.txblkst12                 (txblkst12),                 //   input,   width = 1,           .txblkst12
		.txblkst13                 (txblkst13),                 //   input,   width = 1,           .txblkst13
		.txblkst14                 (txblkst14),                 //   input,   width = 1,           .txblkst14
		.txblkst15                 (txblkst15),                 //   input,   width = 1,           .txblkst15
		.txdataskip8               (txdataskip8),               //   input,   width = 1,           .txdataskip8
		.txdataskip9               (txdataskip9),               //   input,   width = 1,           .txdataskip9
		.txdataskip10              (txdataskip10),              //   input,   width = 1,           .txdataskip10
		.txdataskip11              (txdataskip11),              //   input,   width = 1,           .txdataskip11
		.txdataskip12              (txdataskip12),              //   input,   width = 1,           .txdataskip12
		.txdataskip13              (txdataskip13),              //   input,   width = 1,           .txdataskip13
		.txdataskip14              (txdataskip14),              //   input,   width = 1,           .txdataskip14
		.txdataskip15              (txdataskip15),              //   input,   width = 1,           .txdataskip15
		.rate8                     (rate8),                     //   input,   width = 2,           .rate8
		.rate9                     (rate9),                     //   input,   width = 2,           .rate9
		.rate10                    (rate10),                    //   input,   width = 2,           .rate10
		.rate11                    (rate11),                    //   input,   width = 2,           .rate11
		.rate12                    (rate12),                    //   input,   width = 2,           .rate12
		.rate13                    (rate13),                    //   input,   width = 2,           .rate13
		.rate14                    (rate14),                    //   input,   width = 2,           .rate14
		.rate15                    (rate15),                    //   input,   width = 2,           .rate15
		.test_in                   (test_in),                   //  output,  width = 67,   hip_ctrl.test_in
		.simu_mode_pipe            (simu_mode_pipe),            //  output,   width = 1,           .simu_mode_pipe
		.npor                      (npor),                      //  output,   width = 1,       npor.npor
		.pin_perst                 (pin_perst),                 //  output,   width = 1,           .pin_perst
		.eidleinfersel0            (3'b000),                    // (terminated),                         
		.eidleinfersel1            (3'b000),                    // (terminated),                         
		.eidleinfersel2            (3'b000),                    // (terminated),                         
		.eidleinfersel3            (3'b000),                    // (terminated),                         
		.eidleinfersel4            (3'b000),                    // (terminated),                         
		.eidleinfersel5            (3'b000),                    // (terminated),                         
		.eidleinfersel6            (3'b000),                    // (terminated),                         
		.eidleinfersel7            (3'b000),                    // (terminated),                         
		.eidleinfersel8            (3'b000),                    // (terminated),                         
		.eidleinfersel9            (3'b000),                    // (terminated),                         
		.eidleinfersel10           (3'b000),                    // (terminated),                         
		.eidleinfersel11           (3'b000),                    // (terminated),                         
		.eidleinfersel12           (3'b000),                    // (terminated),                         
		.eidleinfersel13           (3'b000),                    // (terminated),                         
		.eidleinfersel14           (3'b000),                    // (terminated),                         
		.eidleinfersel15           (3'b000)                     // (terminated),                         
	);

endmodule
