// Copyright 2021 Intel Corporation
// SPDX-License-Identifier: MIT

//-----------------------------------------------------------------------------
// Description : List of Tests 
//-----------------------------------------------------------------------------

`ifndef TEST_PKG_SVH
`define TEST_PKG_SVH

//package test_pkg;
//    import uvm_pkg::*;
//    `include "uvm_macros.svh"

    `include "base_test.svh"
    `include "mmio_test.svh"
    `include "he_lpbk_test.svh"
    `include "he_lpbk_long_test.svh"
    `include "he_lpbk_rd_test.svh"
    `include "he_lpbk_wr_test.svh"
    `include "he_lpbk_thruput_test.svh"
    `include "he_lpbk_rd_cont_test.svh"
    `include "he_lpbk_wr_cont_test.svh"
    `include "he_lpbk_thruput_contmode_test.svh"
    `include "he_hssi_csr_test.svh"
    `include "he_mem_lpbk_test.svh"
    `include "he_mem_lpbk_long_test.svh"
    `include "he_mem_wr_test.svh"
    `include "he_mem_rd_test.svh"
    `include "he_mem_thruput_test.svh"
    `include "he_mem_wr_cont_test.svh"
    `include "he_mem_rd_cont_test.svh"
    `include "he_mem_thruput_contmode_test.svh"
    `include "he_mem_cont_test.svh"
    `include "he_hssi_tx_lpbk_test.svh"
    `include "he_hssi_err_test.svh"
    `include "mmio_stress_test.svh"
    `include "he_random_test.svh"
    `include "dfh_walking_test.svh"
    `include "mmio_unimp_test.svh"
    `include "he_lpbk_reqlen1_test.svh"
    `include "he_lpbk_reqlen2_test.svh"
    `include "he_lpbk_reqlen4_test.svh"
    `include "he_lpbk_reqlen8_test.svh"
    `include "he_mem_lpbk_reqlen1_test.svh"
    `include "he_mem_lpbk_reqlen2_test.svh"
    `include "he_mem_lpbk_reqlen4_test.svh"
    `include "he_lpbk_long_rst_test.svh"
    `include "he_mem_lpbk_long_rst_test.svh"
    `include "mmio_stress_nonblocking_test.svh"
    `include "he_lpbk_cont_test.svh"
    `include "fme_csr_test.svh"
    `include "msix_csr_test.svh"
    `include "pmci_csr_test.svh"
    `include "helb_csr_test.svh"
    `include "hemem_csr_test.svh"
    `include "hehssi_csr_test.svh"
    `include "mini_smoke_test.svh"
    `include "mmio_64b_bar_test.svh"
    `include "fme_intr_test.svh"
    `include "flr_reset_test.svh"
    `include "flr_vf0_reset_test.svh"
    `include "flr_vf1_reset_test.svh"
    `include "flr_vf2_reset_test.svh"
    `include "port_gasket_csr_test.svh"
    `include "helb_rd_1cl_test.svh"
    `include "helb_rd_2cl_test.svh"
    `include "helb_rd_4cl_test.svh"
    `include "helb_wr_1cl_test.svh"
    `include "helb_wr_2cl_test.svh"
    `include "helb_wr_4cl_test.svh"
    `include "helb_thruput_1cl_test.svh"
    `include "helb_thruput_2cl_test.svh"
    `include "helb_thruput_4cl_test.svh"
    `include "he_random_long_test.svh"
    `include "hemem_intr_test.svh"
    `include "he_lpbk_port_rst_test.svh"
    `include "fme_hemem_intr_test.svh"
    `include "he_hssi_rx_lpbk_test.svh"
    `include "fme_ras_cat_fat_err_test.svh"
    `include "fme_ras_no_fat_err_test.svh"
     `include "protocol_checker_csr_test.svh"
    `include "MaxTagError_test.svh"
    `include "TxMWrDataPayloadOverrun_test.svh"
    `include "TxMWrInsufficientData_test.svh"
    `include "UnexpMMIORspErr_test.svh"
    `include "malformedtlp_test.svh"
    `include "maxpayloaderror_test.svh"
    `include "MMIOInsufficientData_test.svh"
    `include "MMIOTimedout_test.svh"
    `include "MMIODataPayloadOverrun_test.svh"
    `include "he_mem_user_intr_test.svh"
    `include "he_mem_multi_user_intr_test.svh"

//endpackage : test_pkg

`endif // TEST_PKG_SVH
