// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

`include ".svh"
