`include ".svh"
