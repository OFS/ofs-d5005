// Copyright 2021 Intel Corporation
// SPDX-License-Identifier: MIT

`ifndef RAL_HSSI_SS_CSR
`define RAL_HSSI_SS_CSR

import uvm_pkg::*;

class ral_reg_hssi_ss_csr_HSSI_DFH extends uvm_reg;
	uvm_reg_field FeatureType;
	rand uvm_reg_field Reserved;
	uvm_reg_field EOL;
	uvm_reg_field NextDfhByteOffset;
	uvm_reg_field FeatureRevision;
	uvm_reg_field FeatureId;

	function new(string name = "hssi_ss_csr_HSSI_DFH");
		super.new(name, 64,build_coverage(UVM_NO_COVERAGE));
	endfunction: new
   virtual function void build();
      this.FeatureType = uvm_reg_field::type_id::create("FeatureType",,get_full_name());
      this.FeatureType.configure(this, 4, 60, "RO", 0, 4'h3, 1, 0, 0);
      this.Reserved = uvm_reg_field::type_id::create("Reserved",,get_full_name());
      this.Reserved.configure(this, 19, 41, "WO", 0, 19'h0, 1, 0, 0);
      this.EOL = uvm_reg_field::type_id::create("EOL",,get_full_name());
      this.EOL.configure(this, 1, 40, "RO", 0, 1'h0, 1, 0, 0);
      this.NextDfhByteOffset = uvm_reg_field::type_id::create("NextDfhByteOffset",,get_full_name());
      this.NextDfhByteOffset.configure(this, 24, 16, "RO", 0, 24'h10000, 1, 0, 1);
      this.FeatureRevision = uvm_reg_field::type_id::create("FeatureRevision",,get_full_name());
      this.FeatureRevision.configure(this, 4, 12, "RO", 0, 4'h1, 1, 0, 0);
      this.FeatureId = uvm_reg_field::type_id::create("FeatureId",,get_full_name());
      this.FeatureId.configure(this, 4, 12, "RO", 0, 4'h1, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_hssi_ss_csr_HSSI_DFH)

endclass : ral_reg_hssi_ss_csr_HSSI_DFH


class ral_reg_hssi_ss_csr_HSSI_CAPABILITY extends uvm_reg;
	rand uvm_reg_field Reserved;
	uvm_reg_field NumQSFPInterfaces;
	uvm_reg_field num_channels;
	uvm_reg_field Num_channels_CSR_interface;
	uvm_reg_field Num_CSR_interface;

	function new(string name = "hssi_ss_csr_HSSI_CAPABILITY");
		super.new(name, 64,build_coverage(UVM_NO_COVERAGE));
	endfunction: new
   virtual function void build();
      this.Reserved = uvm_reg_field::type_id::create("Reserved",,get_full_name());
      this.Reserved.configure(this, 20, 44, "WO", 0, 20'h0, 1, 0, 0);
      this.NumQSFPInterfaces = uvm_reg_field::type_id::create("NumQSFPInterfaces",,get_full_name());
      this.NumQSFPInterfaces.configure(this, 4, 40, "RO", 0, 4'h0, 1, 0, 0);
      this.num_channels = uvm_reg_field::type_id::create("num_channels",,get_full_name());
      this.num_channels.configure(this, 4, 36, "RO", 0, 4'h0, 1, 0, 0);
      this.Num_channels_CSR_interface = uvm_reg_field::type_id::create("Num_channels_CSR_interface",,get_full_name());
      this.Num_channels_CSR_interface.configure(this, 4, 32, "RO", 0, 4'h2, 1, 0, 0);
      this.Num_CSR_interface = uvm_reg_field::type_id::create("Num_CSR_interface",,get_full_name());
      this.Num_CSR_interface.configure(this, 4, 28, "RO", 0, 4'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_hssi_ss_csr_HSSI_CAPABILITY)

endclass : ral_reg_hssi_ss_csr_HSSI_CAPABILITY


class ral_reg_hssi_ss_csr_HSSI_CTRL extends uvm_reg;
	rand uvm_reg_field Reserved;

	function new(string name = "hssi_ss_csr_HSSI_CTRL");
		super.new(name, 64,build_coverage(UVM_NO_COVERAGE));
	endfunction: new
   virtual function void build();
      this.Reserved = uvm_reg_field::type_id::create("Reserved",,get_full_name());
      this.Reserved.configure(this, 36, 28, "WO", 0, 36'h000000000, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_hssi_ss_csr_HSSI_CTRL)

endclass : ral_reg_hssi_ss_csr_HSSI_CTRL


class ral_reg_hssi_ss_csr_HSSI_STAT0 extends uvm_reg;
	uvm_reg_field Chan3RxReady;
	uvm_reg_field Chan3TxReady;
	uvm_reg_field Chan3RxIsLockedToRef;
	uvm_reg_field Chan3RxIsLockedToData;
	uvm_reg_field EChan3RxCalBusy;
	uvm_reg_field Chan3TxCalBusy;
	uvm_reg_field Chan3RxTransferReady;
	uvm_reg_field Chan3TxTransferReady;
	uvm_reg_field Chan3RxFifoReady;
	uvm_reg_field Chan3TxFifoReady;
	uvm_reg_field Chan3RxDigitalResetTimeout;
	uvm_reg_field Chan3TxDigitalResetTimeout;
	uvm_reg_field Chan3RxDigitalResetStat;
	uvm_reg_field Chan3RxAnalogResetStat;
	uvm_reg_field Chan3TxDigitalResetStat;
	uvm_reg_field Chan3TxAnalogResetStat;
	uvm_reg_field Chan2RxReady;
	uvm_reg_field Chan2TxReady;
	uvm_reg_field Chan2RxIsLockedToRef;
	uvm_reg_field Chan2RxIsLockedToData;
	uvm_reg_field Chan2RxCalBusy;
	uvm_reg_field Chan2TxCalBusy;
	uvm_reg_field Chan2RxTransferReady;
	uvm_reg_field Chan2TxTransferReady;
	uvm_reg_field Chan2RxFifoReady;
	uvm_reg_field Chan2TxFifoReady;
	uvm_reg_field Chan2RxDigitalResetTimeout;
	uvm_reg_field Chan2TxDigitalResetTimeout;
	uvm_reg_field Chan2RxDigitalResetStat;
	uvm_reg_field Chan2RxAnalogResetStat;
	uvm_reg_field Chan2TxDigitalResetStat;
	uvm_reg_field Chan2TxAnalogResetStat;
	uvm_reg_field Chan1RxReady;
	uvm_reg_field Chan1TxReady;
	uvm_reg_field Chan1RxIsLockedToRef;
	uvm_reg_field Chan1RxIsLockedToData;
	uvm_reg_field Chan1RxCalBusy;
	uvm_reg_field Chan1TxCalBusy;
	uvm_reg_field Chan1RxTransferReady;
	uvm_reg_field Chan1TxTransferReady;
	uvm_reg_field Chan1RxFifoReady;
	uvm_reg_field Chan1TxFifoReady;
	uvm_reg_field Chan1RxDigitalResetTimeout;
	uvm_reg_field Chan1TxDigitalResetTimeout;
	uvm_reg_field Chan1RxDigitalResetStat;
	uvm_reg_field Chan1RxAnalogResetStat;
	uvm_reg_field Chan1TxDigitalResetStat;
	uvm_reg_field Chan1TxAnalogResetStat;
	uvm_reg_field Chan0RxReady;
	uvm_reg_field Chan0TxReady;
	uvm_reg_field Chan0RxIsLockedToRef;
	uvm_reg_field Chan0RxIsLockedToData;
	uvm_reg_field Chan0RxCalBusy;
	uvm_reg_field Chan0TxCalBusy;
	uvm_reg_field Chan0RxTransferReady;
	uvm_reg_field Chan0TxTransferReady;
	uvm_reg_field Chan0RxFifoReady;
	uvm_reg_field Chan0TxFifoReady;
	uvm_reg_field Chan0RxDigitalResetTimeout;
	uvm_reg_field Chan0TxDigitalResetTimeout;
	uvm_reg_field Chan0RxDigitalResetStat;
	uvm_reg_field Chan0RxAnalogResetStat;
	uvm_reg_field Chan0TxDigitalResetStat;
	uvm_reg_field Chan0TxAnalogResetStat;

	function new(string name = "hssi_ss_csr_HSSI_STAT0");
		super.new(name, 64,build_coverage(UVM_NO_COVERAGE));
	endfunction: new
   virtual function void build();
      this.Chan3RxReady = uvm_reg_field::type_id::create("Chan3RxReady",,get_full_name());
      this.Chan3RxReady.configure(this, 1, 63, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3TxReady = uvm_reg_field::type_id::create("Chan3TxReady",,get_full_name());
      this.Chan3TxReady.configure(this, 1, 62, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3RxIsLockedToRef = uvm_reg_field::type_id::create("Chan3RxIsLockedToRef",,get_full_name());
      this.Chan3RxIsLockedToRef.configure(this, 1, 61, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3RxIsLockedToData = uvm_reg_field::type_id::create("Chan3RxIsLockedToData",,get_full_name());
      this.Chan3RxIsLockedToData.configure(this, 1, 60, "RO", 0, 1'h0, 1, 0, 0);
      this.EChan3RxCalBusy = uvm_reg_field::type_id::create("EChan3RxCalBusy",,get_full_name());
      this.EChan3RxCalBusy.configure(this, 1, 59, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3TxCalBusy = uvm_reg_field::type_id::create("Chan3TxCalBusy",,get_full_name());
      this.Chan3TxCalBusy.configure(this, 1, 58, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3RxTransferReady = uvm_reg_field::type_id::create("Chan3RxTransferReady",,get_full_name());
      this.Chan3RxTransferReady.configure(this, 1, 57, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3TxTransferReady = uvm_reg_field::type_id::create("Chan3TxTransferReady",,get_full_name());
      this.Chan3TxTransferReady.configure(this, 1, 56, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3RxFifoReady = uvm_reg_field::type_id::create("Chan3RxFifoReady",,get_full_name());
      this.Chan3RxFifoReady.configure(this, 1, 55, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3TxFifoReady = uvm_reg_field::type_id::create("Chan3TxFifoReady",,get_full_name());
      this.Chan3TxFifoReady.configure(this, 1, 54, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3RxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan3RxDigitalResetTimeout",,get_full_name());
      this.Chan3RxDigitalResetTimeout.configure(this, 1, 53, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3TxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan3TxDigitalResetTimeout",,get_full_name());
      this.Chan3TxDigitalResetTimeout.configure(this, 1, 52, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3RxDigitalResetStat = uvm_reg_field::type_id::create("Chan3RxDigitalResetStat",,get_full_name());
      this.Chan3RxDigitalResetStat.configure(this, 1, 51, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3RxAnalogResetStat = uvm_reg_field::type_id::create("Chan3RxAnalogResetStat",,get_full_name());
      this.Chan3RxAnalogResetStat.configure(this, 1, 50, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3TxDigitalResetStat = uvm_reg_field::type_id::create("Chan3TxDigitalResetStat",,get_full_name());
      this.Chan3TxDigitalResetStat.configure(this, 1, 49, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan3TxAnalogResetStat = uvm_reg_field::type_id::create("Chan3TxAnalogResetStat",,get_full_name());
      this.Chan3TxAnalogResetStat.configure(this, 1, 48, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxReady = uvm_reg_field::type_id::create("Chan2RxReady",,get_full_name());
      this.Chan2RxReady.configure(this, 1, 47, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2TxReady = uvm_reg_field::type_id::create("Chan2TxReady",,get_full_name());
      this.Chan2TxReady.configure(this, 1, 46, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxIsLockedToRef = uvm_reg_field::type_id::create("Chan2RxIsLockedToRef",,get_full_name());
      this.Chan2RxIsLockedToRef.configure(this, 1, 45, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxIsLockedToData = uvm_reg_field::type_id::create("Chan2RxIsLockedToData",,get_full_name());
      this.Chan2RxIsLockedToData.configure(this, 1, 44, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxCalBusy = uvm_reg_field::type_id::create("Chan2RxCalBusy",,get_full_name());
      this.Chan2RxCalBusy.configure(this, 1, 43, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2TxCalBusy = uvm_reg_field::type_id::create("Chan2TxCalBusy",,get_full_name());
      this.Chan2TxCalBusy.configure(this, 1, 42, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxTransferReady = uvm_reg_field::type_id::create("Chan2RxTransferReady",,get_full_name());
      this.Chan2RxTransferReady.configure(this, 1, 41, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2TxTransferReady = uvm_reg_field::type_id::create("Chan2TxTransferReady",,get_full_name());
      this.Chan2TxTransferReady.configure(this, 1, 40, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxFifoReady = uvm_reg_field::type_id::create("Chan2RxFifoReady",,get_full_name());
      this.Chan2RxFifoReady.configure(this, 1, 39, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2TxFifoReady = uvm_reg_field::type_id::create("Chan2TxFifoReady",,get_full_name());
      this.Chan2TxFifoReady.configure(this, 1, 38, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan2RxDigitalResetTimeout",,get_full_name());
      this.Chan2RxDigitalResetTimeout.configure(this, 1, 37, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2TxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan2TxDigitalResetTimeout",,get_full_name());
      this.Chan2TxDigitalResetTimeout.configure(this, 1, 36, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxDigitalResetStat = uvm_reg_field::type_id::create("Chan2RxDigitalResetStat",,get_full_name());
      this.Chan2RxDigitalResetStat.configure(this, 1, 35, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2RxAnalogResetStat = uvm_reg_field::type_id::create("Chan2RxAnalogResetStat",,get_full_name());
      this.Chan2RxAnalogResetStat.configure(this, 1, 34, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2TxDigitalResetStat = uvm_reg_field::type_id::create("Chan2TxDigitalResetStat",,get_full_name());
      this.Chan2TxDigitalResetStat.configure(this, 1, 33, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan2TxAnalogResetStat = uvm_reg_field::type_id::create("Chan2TxAnalogResetStat",,get_full_name());
      this.Chan2TxAnalogResetStat.configure(this, 1, 32, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxReady = uvm_reg_field::type_id::create("Chan1RxReady",,get_full_name());
      this.Chan1RxReady.configure(this, 1, 31, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1TxReady = uvm_reg_field::type_id::create("Chan1TxReady",,get_full_name());
      this.Chan1TxReady.configure(this, 1, 30, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxIsLockedToRef = uvm_reg_field::type_id::create("Chan1RxIsLockedToRef",,get_full_name());
      this.Chan1RxIsLockedToRef.configure(this, 1, 29, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxIsLockedToData = uvm_reg_field::type_id::create("Chan1RxIsLockedToData",,get_full_name());
      this.Chan1RxIsLockedToData.configure(this, 1, 28, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxCalBusy = uvm_reg_field::type_id::create("Chan1RxCalBusy",,get_full_name());
      this.Chan1RxCalBusy.configure(this, 1, 27, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1TxCalBusy = uvm_reg_field::type_id::create("Chan1TxCalBusy",,get_full_name());
      this.Chan1TxCalBusy.configure(this, 1, 26, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxTransferReady = uvm_reg_field::type_id::create("Chan1RxTransferReady",,get_full_name());
      this.Chan1RxTransferReady.configure(this, 1, 25, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1TxTransferReady = uvm_reg_field::type_id::create("Chan1TxTransferReady",,get_full_name());
      this.Chan1TxTransferReady.configure(this, 1, 24, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxFifoReady = uvm_reg_field::type_id::create("Chan1RxFifoReady",,get_full_name());
      this.Chan1RxFifoReady.configure(this, 1, 23, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1TxFifoReady = uvm_reg_field::type_id::create("Chan1TxFifoReady",,get_full_name());
      this.Chan1TxFifoReady.configure(this, 1, 22, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan1RxDigitalResetTimeout",,get_full_name());
      this.Chan1RxDigitalResetTimeout.configure(this, 1, 21, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1TxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan1TxDigitalResetTimeout",,get_full_name());
      this.Chan1TxDigitalResetTimeout.configure(this, 1, 20, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxDigitalResetStat = uvm_reg_field::type_id::create("Chan1RxDigitalResetStat",,get_full_name());
      this.Chan1RxDigitalResetStat.configure(this, 1, 19, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1RxAnalogResetStat = uvm_reg_field::type_id::create("Chan1RxAnalogResetStat",,get_full_name());
      this.Chan1RxAnalogResetStat.configure(this, 1, 18, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1TxDigitalResetStat = uvm_reg_field::type_id::create("Chan1TxDigitalResetStat",,get_full_name());
      this.Chan1TxDigitalResetStat.configure(this, 1, 17, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1TxAnalogResetStat = uvm_reg_field::type_id::create("Chan1TxAnalogResetStat",,get_full_name());
      this.Chan1TxAnalogResetStat.configure(this, 1, 16, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxReady = uvm_reg_field::type_id::create("Chan0RxReady",,get_full_name());
      this.Chan0RxReady.configure(this, 1, 15, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0TxReady = uvm_reg_field::type_id::create("Chan0TxReady",,get_full_name());
      this.Chan0TxReady.configure(this, 1, 14, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxIsLockedToRef = uvm_reg_field::type_id::create("Chan0RxIsLockedToRef",,get_full_name());
      this.Chan0RxIsLockedToRef.configure(this, 1, 13, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxIsLockedToData = uvm_reg_field::type_id::create("Chan0RxIsLockedToData",,get_full_name());
      this.Chan0RxIsLockedToData.configure(this, 1, 12, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxCalBusy = uvm_reg_field::type_id::create("Chan0RxCalBusy",,get_full_name());
      this.Chan0RxCalBusy.configure(this, 1, 11, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0TxCalBusy = uvm_reg_field::type_id::create("Chan0TxCalBusy",,get_full_name());
      this.Chan0TxCalBusy.configure(this, 1, 10, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxTransferReady = uvm_reg_field::type_id::create("Chan0RxTransferReady",,get_full_name());
      this.Chan0RxTransferReady.configure(this, 1, 9, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0TxTransferReady = uvm_reg_field::type_id::create("Chan0TxTransferReady",,get_full_name());
      this.Chan0TxTransferReady.configure(this, 1, 8, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxFifoReady = uvm_reg_field::type_id::create("Chan0RxFifoReady",,get_full_name());
      this.Chan0RxFifoReady.configure(this, 1, 7, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0TxFifoReady = uvm_reg_field::type_id::create("Chan0TxFifoReady",,get_full_name());
      this.Chan0TxFifoReady.configure(this, 1, 6, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan0RxDigitalResetTimeout",,get_full_name());
      this.Chan0RxDigitalResetTimeout.configure(this, 1, 5, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0TxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan0TxDigitalResetTimeout",,get_full_name());
      this.Chan0TxDigitalResetTimeout.configure(this, 1, 4, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxDigitalResetStat = uvm_reg_field::type_id::create("Chan0RxDigitalResetStat",,get_full_name());
      this.Chan0RxDigitalResetStat.configure(this, 1, 3, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0RxAnalogResetStat = uvm_reg_field::type_id::create("Chan0RxAnalogResetStat",,get_full_name());
      this.Chan0RxAnalogResetStat.configure(this, 1, 2, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0TxDigitalResetStat = uvm_reg_field::type_id::create("Chan0TxDigitalResetStat",,get_full_name());
      this.Chan0TxDigitalResetStat.configure(this, 1, 1, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan0TxAnalogResetStat = uvm_reg_field::type_id::create("Chan0TxAnalogResetStat",,get_full_name());
      this.Chan0TxAnalogResetStat.configure(this, 1, 0, "RO", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_hssi_ss_csr_HSSI_STAT0)

endclass : ral_reg_hssi_ss_csr_HSSI_STAT0


class ral_reg_hssi_ss_csr_HSSI_STAT1 extends uvm_reg;
	uvm_reg_field Chan7RxReady;
	uvm_reg_field Chan7TxReady;
	uvm_reg_field Chan7RxIsLockedToRef;
	uvm_reg_field Chan7RxIsLockedToData;
	uvm_reg_field EChan7RxCalBusy;
	uvm_reg_field Chan7TxCalBusy;
	uvm_reg_field Chan7RxTransferReady;
	uvm_reg_field Chan7TxTransferReady;
	uvm_reg_field Chan7RxFifoReady;
	uvm_reg_field Chan7TxFifoReady;
	uvm_reg_field Chan7RxDigitalResetTimeout;
	uvm_reg_field Chan7TxDigitalResetTimeout;
	uvm_reg_field Chan7RxDigitalResetStat;
	uvm_reg_field Chan7RxAnalogResetStat;
	uvm_reg_field Chan7TxDigitalResetStat;
	uvm_reg_field Chan7TxAnalogResetStat;
	uvm_reg_field Chan6RxReady;
	uvm_reg_field Chan6TxReady;
	uvm_reg_field Chan6RxIsLockedToRef;
	uvm_reg_field Chan6RxIsLockedToData;
	uvm_reg_field Chan6RxCalBusy;
	uvm_reg_field Chan6TxCalBusy;
	uvm_reg_field Chan6RxTransferReady;
	uvm_reg_field Chan6TxTransferReady;
	uvm_reg_field Chan6RxFifoReady;
	uvm_reg_field Chan6TxFifoReady;
	uvm_reg_field Chan6RxDigitalResetTimeout;
	uvm_reg_field Chan6TxDigitalResetTimeout;
	uvm_reg_field Chan6RxDigitalResetStat;
	uvm_reg_field Chan6RxAnalogResetStat;
	uvm_reg_field Chan6TxDigitalResetStat;
	uvm_reg_field Chan6TxAnalogResetStat;
	uvm_reg_field Chan5RxReady;
	uvm_reg_field Chan5TxReady;
	uvm_reg_field Chan5RxIsLockedToRef;
	uvm_reg_field Chan5RxIsLockedToData;
	uvm_reg_field Chan5RxCalBusy;
	uvm_reg_field Chan1TxCalBusy;
	uvm_reg_field Chan5RxTransferReady;
	uvm_reg_field Chan5TxTransferReady;
	uvm_reg_field Chan5RxFifoReady;
	uvm_reg_field Chan5TxFifoReady;
	uvm_reg_field Chan5RxDigitalResetTimeout;
	uvm_reg_field Chan5TxDigitalResetTimeout;
	uvm_reg_field Chan5RxDigitalResetStat;
	uvm_reg_field Chan5RxAnalogResetStat;
	uvm_reg_field Chan5TxDigitalResetStat;
	uvm_reg_field Chan5TxAnalogResetStat;
	uvm_reg_field Chan4RxReady;
	uvm_reg_field Chan4TxReady;
	uvm_reg_field Chan4RxIsLockedToRef;
	uvm_reg_field Chan4RxIsLockedToData;
	uvm_reg_field Chan4RxCalBusy;
	uvm_reg_field Chan4TxCalBusy;
	uvm_reg_field Chan4RxTransferReady;
	uvm_reg_field Chan4TxTransferReady;
	uvm_reg_field Chan4RxFifoReady;
	uvm_reg_field Chan4TxFifoReady;
	uvm_reg_field Chan4RxDigitalResetTimeout;
	uvm_reg_field Chan4TxDigitalResetTimeout;
	uvm_reg_field Chan4RxDigitalResetStat;
	uvm_reg_field Chan4RxAnalogResetStat;
	uvm_reg_field Chan4TxDigitalResetStat;
	uvm_reg_field Chan4TxAnalogResetStat;

	function new(string name = "hssi_ss_csr_HSSI_STAT1");
		super.new(name, 64,build_coverage(UVM_NO_COVERAGE));
	endfunction: new
   virtual function void build();
      this.Chan7RxReady = uvm_reg_field::type_id::create("Chan7RxReady",,get_full_name());
      this.Chan7RxReady.configure(this, 1, 63, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7TxReady = uvm_reg_field::type_id::create("Chan7TxReady",,get_full_name());
      this.Chan7TxReady.configure(this, 1, 62, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7RxIsLockedToRef = uvm_reg_field::type_id::create("Chan7RxIsLockedToRef",,get_full_name());
      this.Chan7RxIsLockedToRef.configure(this, 1, 61, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7RxIsLockedToData = uvm_reg_field::type_id::create("Chan7RxIsLockedToData",,get_full_name());
      this.Chan7RxIsLockedToData.configure(this, 1, 60, "RO", 0, 1'h0, 1, 0, 0);
      this.EChan7RxCalBusy = uvm_reg_field::type_id::create("EChan7RxCalBusy",,get_full_name());
      this.EChan7RxCalBusy.configure(this, 1, 59, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7TxCalBusy = uvm_reg_field::type_id::create("Chan7TxCalBusy",,get_full_name());
      this.Chan7TxCalBusy.configure(this, 1, 58, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7RxTransferReady = uvm_reg_field::type_id::create("Chan7RxTransferReady",,get_full_name());
      this.Chan7RxTransferReady.configure(this, 1, 57, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7TxTransferReady = uvm_reg_field::type_id::create("Chan7TxTransferReady",,get_full_name());
      this.Chan7TxTransferReady.configure(this, 1, 56, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7RxFifoReady = uvm_reg_field::type_id::create("Chan7RxFifoReady",,get_full_name());
      this.Chan7RxFifoReady.configure(this, 1, 55, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7TxFifoReady = uvm_reg_field::type_id::create("Chan7TxFifoReady",,get_full_name());
      this.Chan7TxFifoReady.configure(this, 1, 54, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7RxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan7RxDigitalResetTimeout",,get_full_name());
      this.Chan7RxDigitalResetTimeout.configure(this, 1, 53, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7TxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan7TxDigitalResetTimeout",,get_full_name());
      this.Chan7TxDigitalResetTimeout.configure(this, 1, 52, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7RxDigitalResetStat = uvm_reg_field::type_id::create("Chan7RxDigitalResetStat",,get_full_name());
      this.Chan7RxDigitalResetStat.configure(this, 1, 51, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7RxAnalogResetStat = uvm_reg_field::type_id::create("Chan7RxAnalogResetStat",,get_full_name());
      this.Chan7RxAnalogResetStat.configure(this, 1, 50, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7TxDigitalResetStat = uvm_reg_field::type_id::create("Chan7TxDigitalResetStat",,get_full_name());
      this.Chan7TxDigitalResetStat.configure(this, 1, 49, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan7TxAnalogResetStat = uvm_reg_field::type_id::create("Chan7TxAnalogResetStat",,get_full_name());
      this.Chan7TxAnalogResetStat.configure(this, 1, 48, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxReady = uvm_reg_field::type_id::create("Chan6RxReady",,get_full_name());
      this.Chan6RxReady.configure(this, 1, 47, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6TxReady = uvm_reg_field::type_id::create("Chan6TxReady",,get_full_name());
      this.Chan6TxReady.configure(this, 1, 46, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxIsLockedToRef = uvm_reg_field::type_id::create("Chan6RxIsLockedToRef",,get_full_name());
      this.Chan6RxIsLockedToRef.configure(this, 1, 45, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxIsLockedToData = uvm_reg_field::type_id::create("Chan6RxIsLockedToData",,get_full_name());
      this.Chan6RxIsLockedToData.configure(this, 1, 44, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxCalBusy = uvm_reg_field::type_id::create("Chan6RxCalBusy",,get_full_name());
      this.Chan6RxCalBusy.configure(this, 1, 43, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6TxCalBusy = uvm_reg_field::type_id::create("Chan6TxCalBusy",,get_full_name());
      this.Chan6TxCalBusy.configure(this, 1, 42, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxTransferReady = uvm_reg_field::type_id::create("Chan6RxTransferReady",,get_full_name());
      this.Chan6RxTransferReady.configure(this, 1, 41, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6TxTransferReady = uvm_reg_field::type_id::create("Chan6TxTransferReady",,get_full_name());
      this.Chan6TxTransferReady.configure(this, 1, 40, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxFifoReady = uvm_reg_field::type_id::create("Chan6RxFifoReady",,get_full_name());
      this.Chan6RxFifoReady.configure(this, 1, 39, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6TxFifoReady = uvm_reg_field::type_id::create("Chan6TxFifoReady",,get_full_name());
      this.Chan6TxFifoReady.configure(this, 1, 38, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan6RxDigitalResetTimeout",,get_full_name());
      this.Chan6RxDigitalResetTimeout.configure(this, 1, 37, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6TxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan6TxDigitalResetTimeout",,get_full_name());
      this.Chan6TxDigitalResetTimeout.configure(this, 1, 36, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxDigitalResetStat = uvm_reg_field::type_id::create("Chan6RxDigitalResetStat",,get_full_name());
      this.Chan6RxDigitalResetStat.configure(this, 1, 35, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6RxAnalogResetStat = uvm_reg_field::type_id::create("Chan6RxAnalogResetStat",,get_full_name());
      this.Chan6RxAnalogResetStat.configure(this, 1, 34, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6TxDigitalResetStat = uvm_reg_field::type_id::create("Chan6TxDigitalResetStat",,get_full_name());
      this.Chan6TxDigitalResetStat.configure(this, 1, 33, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan6TxAnalogResetStat = uvm_reg_field::type_id::create("Chan6TxAnalogResetStat",,get_full_name());
      this.Chan6TxAnalogResetStat.configure(this, 1, 32, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxReady = uvm_reg_field::type_id::create("Chan5RxReady",,get_full_name());
      this.Chan5RxReady.configure(this, 1, 31, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5TxReady = uvm_reg_field::type_id::create("Chan5TxReady",,get_full_name());
      this.Chan5TxReady.configure(this, 1, 30, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxIsLockedToRef = uvm_reg_field::type_id::create("Chan5RxIsLockedToRef",,get_full_name());
      this.Chan5RxIsLockedToRef.configure(this, 1, 29, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxIsLockedToData = uvm_reg_field::type_id::create("Chan5RxIsLockedToData",,get_full_name());
      this.Chan5RxIsLockedToData.configure(this, 1, 28, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxCalBusy = uvm_reg_field::type_id::create("Chan5RxCalBusy",,get_full_name());
      this.Chan5RxCalBusy.configure(this, 1, 27, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan1TxCalBusy = uvm_reg_field::type_id::create("Chan1TxCalBusy",,get_full_name());
      this.Chan1TxCalBusy.configure(this, 1, 26, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxTransferReady = uvm_reg_field::type_id::create("Chan5RxTransferReady",,get_full_name());
      this.Chan5RxTransferReady.configure(this, 1, 25, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5TxTransferReady = uvm_reg_field::type_id::create("Chan5TxTransferReady",,get_full_name());
      this.Chan5TxTransferReady.configure(this, 1, 24, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxFifoReady = uvm_reg_field::type_id::create("Chan5RxFifoReady",,get_full_name());
      this.Chan5RxFifoReady.configure(this, 1, 23, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5TxFifoReady = uvm_reg_field::type_id::create("Chan5TxFifoReady",,get_full_name());
      this.Chan5TxFifoReady.configure(this, 1, 22, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan5RxDigitalResetTimeout",,get_full_name());
      this.Chan5RxDigitalResetTimeout.configure(this, 1, 21, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5TxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan5TxDigitalResetTimeout",,get_full_name());
      this.Chan5TxDigitalResetTimeout.configure(this, 1, 20, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxDigitalResetStat = uvm_reg_field::type_id::create("Chan5RxDigitalResetStat",,get_full_name());
      this.Chan5RxDigitalResetStat.configure(this, 1, 19, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5RxAnalogResetStat = uvm_reg_field::type_id::create("Chan5RxAnalogResetStat",,get_full_name());
      this.Chan5RxAnalogResetStat.configure(this, 1, 18, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5TxDigitalResetStat = uvm_reg_field::type_id::create("Chan5TxDigitalResetStat",,get_full_name());
      this.Chan5TxDigitalResetStat.configure(this, 1, 17, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan5TxAnalogResetStat = uvm_reg_field::type_id::create("Chan5TxAnalogResetStat",,get_full_name());
      this.Chan5TxAnalogResetStat.configure(this, 1, 16, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxReady = uvm_reg_field::type_id::create("Chan4RxReady",,get_full_name());
      this.Chan4RxReady.configure(this, 1, 15, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4TxReady = uvm_reg_field::type_id::create("Chan4TxReady",,get_full_name());
      this.Chan4TxReady.configure(this, 1, 14, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxIsLockedToRef = uvm_reg_field::type_id::create("Chan4RxIsLockedToRef",,get_full_name());
      this.Chan4RxIsLockedToRef.configure(this, 1, 13, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxIsLockedToData = uvm_reg_field::type_id::create("Chan4RxIsLockedToData",,get_full_name());
      this.Chan4RxIsLockedToData.configure(this, 1, 12, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxCalBusy = uvm_reg_field::type_id::create("Chan4RxCalBusy",,get_full_name());
      this.Chan4RxCalBusy.configure(this, 1, 11, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4TxCalBusy = uvm_reg_field::type_id::create("Chan4TxCalBusy",,get_full_name());
      this.Chan4TxCalBusy.configure(this, 1, 10, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxTransferReady = uvm_reg_field::type_id::create("Chan4RxTransferReady",,get_full_name());
      this.Chan4RxTransferReady.configure(this, 1, 9, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4TxTransferReady = uvm_reg_field::type_id::create("Chan4TxTransferReady",,get_full_name());
      this.Chan4TxTransferReady.configure(this, 1, 8, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxFifoReady = uvm_reg_field::type_id::create("Chan4RxFifoReady",,get_full_name());
      this.Chan4RxFifoReady.configure(this, 1, 7, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4TxFifoReady = uvm_reg_field::type_id::create("Chan4TxFifoReady",,get_full_name());
      this.Chan4TxFifoReady.configure(this, 1, 6, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan4RxDigitalResetTimeout",,get_full_name());
      this.Chan4RxDigitalResetTimeout.configure(this, 1, 5, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4TxDigitalResetTimeout = uvm_reg_field::type_id::create("Chan4TxDigitalResetTimeout",,get_full_name());
      this.Chan4TxDigitalResetTimeout.configure(this, 1, 4, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxDigitalResetStat = uvm_reg_field::type_id::create("Chan4RxDigitalResetStat",,get_full_name());
      this.Chan4RxDigitalResetStat.configure(this, 1, 3, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4RxAnalogResetStat = uvm_reg_field::type_id::create("Chan4RxAnalogResetStat",,get_full_name());
      this.Chan4RxAnalogResetStat.configure(this, 1, 2, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4TxDigitalResetStat = uvm_reg_field::type_id::create("Chan4TxDigitalResetStat",,get_full_name());
      this.Chan4TxDigitalResetStat.configure(this, 1, 1, "RO", 0, 1'h0, 1, 0, 0);
      this.Chan4TxAnalogResetStat = uvm_reg_field::type_id::create("Chan4TxAnalogResetStat",,get_full_name());
      this.Chan4TxAnalogResetStat.configure(this, 1, 0, "RO", 0, 1'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_hssi_ss_csr_HSSI_STAT1)

endclass : ral_reg_hssi_ss_csr_HSSI_STAT1


class ral_reg_hssi_ss_csr_HSSI_RCFG_CMD0 extends uvm_reg;
	rand uvm_reg_field Reserved;
	rand uvm_reg_field XcvrRcfgAddr;
	rand uvm_reg_field Reserved_1;
	uvm_reg_field XcvrRcfgAck;
	rand uvm_reg_field XcvrRcfgCmdStatus;

	function new(string name = "hssi_ss_csr_HSSI_RCFG_CMD0");
		super.new(name, 64,build_coverage(UVM_NO_COVERAGE));
	endfunction: new
   virtual function void build();
      this.Reserved = uvm_reg_field::type_id::create("Reserved",,get_full_name());
      this.Reserved.configure(this, 12, 52, "WO", 0, 12'h0, 1, 0, 0);
      this.XcvrRcfgAddr = uvm_reg_field::type_id::create("XcvrRcfgAddr",,get_full_name());
      this.XcvrRcfgAddr.configure(this, 20, 32, "RW", 0, 20'h0, 1, 0, 0);
      this.Reserved_1 = uvm_reg_field::type_id::create("Reserved_1",,get_full_name());
      this.Reserved_1.configure(this, 29, 3, "WO", 0, 29'h0, 1, 0, 0);
      this.XcvrRcfgAck = uvm_reg_field::type_id::create("XcvrRcfgAck",,get_full_name());
      this.XcvrRcfgAck.configure(this, 1, 2, "RO", 0, 1'h0, 1, 0, 0);
      this.XcvrRcfgCmdStatus = uvm_reg_field::type_id::create("XcvrRcfgCmdStatus",,get_full_name());
      this.XcvrRcfgCmdStatus.configure(this, 2, 0, "RW", 0, 2'h0, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_hssi_ss_csr_HSSI_RCFG_CMD0)

endclass : ral_reg_hssi_ss_csr_HSSI_RCFG_CMD0


class ral_reg_hssi_ss_csr_HSSI_RCFG_DATA0 extends uvm_reg;
	rand uvm_reg_field XcvrRcfgWrData;
	uvm_reg_field XcvrRcfgRdData;

	function new(string name = "hssi_ss_csr_HSSI_RCFG_DATA0");
		super.new(name, 64,build_coverage(UVM_NO_COVERAGE));
	endfunction: new
   virtual function void build();
      this.XcvrRcfgWrData = uvm_reg_field::type_id::create("XcvrRcfgWrData",,get_full_name());
      this.XcvrRcfgWrData.configure(this, 32, 32, "RW", 0, 32'h0, 1, 0, 1);
      this.XcvrRcfgRdData = uvm_reg_field::type_id::create("XcvrRcfgRdData",,get_full_name());
      this.XcvrRcfgRdData.configure(this, 32, 0, "RO", 0, 32'h0, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_hssi_ss_csr_HSSI_RCFG_DATA0)

endclass : ral_reg_hssi_ss_csr_HSSI_RCFG_DATA0


class ral_reg_hssi_ss_csr_HSSI_SCRATCHPAD extends uvm_reg;
	rand uvm_reg_field Scrathpad;

	function new(string name = "hssi_ss_csr_HSSI_SCRATCHPAD");
		super.new(name, 64,build_coverage(UVM_NO_COVERAGE));
	endfunction: new
   virtual function void build();
      this.Scrathpad = uvm_reg_field::type_id::create("Scrathpad",,get_full_name());
      this.Scrathpad.configure(this, 64, 0, "RW", 0, 64'h000000000, 1, 0, 1);
   endfunction: build

	`uvm_object_utils(ral_reg_hssi_ss_csr_HSSI_SCRATCHPAD)

endclass : ral_reg_hssi_ss_csr_HSSI_SCRATCHPAD


class ral_block_hssi_ss_csr extends uvm_reg_block;
	rand ral_reg_hssi_ss_csr_HSSI_DFH HSSI_DFH;
	rand ral_reg_hssi_ss_csr_HSSI_CAPABILITY HSSI_CAPABILITY;
	rand ral_reg_hssi_ss_csr_HSSI_CTRL HSSI_CTRL;
	rand ral_reg_hssi_ss_csr_HSSI_STAT0 HSSI_STAT0;
	rand ral_reg_hssi_ss_csr_HSSI_STAT1 HSSI_STAT1;
	rand ral_reg_hssi_ss_csr_HSSI_RCFG_CMD0 HSSI_RCFG_CMD0;
	rand ral_reg_hssi_ss_csr_HSSI_RCFG_DATA0 HSSI_RCFG_DATA0;
	rand ral_reg_hssi_ss_csr_HSSI_SCRATCHPAD HSSI_SCRATCHPAD;
	uvm_reg_field HSSI_DFH_FeatureType;
	uvm_reg_field FeatureType;
	rand uvm_reg_field HSSI_DFH_Reserved;
	uvm_reg_field HSSI_DFH_EOL;
	uvm_reg_field EOL;
	uvm_reg_field HSSI_DFH_NextDfhByteOffset;
	uvm_reg_field NextDfhByteOffset;
	uvm_reg_field HSSI_DFH_FeatureRevision;
	uvm_reg_field FeatureRevision;
	uvm_reg_field HSSI_DFH_FeatureId;
	uvm_reg_field FeatureId;
	rand uvm_reg_field HSSI_CAPABILITY_Reserved;
	uvm_reg_field HSSI_CAPABILITY_NumQSFPInterfaces;
	uvm_reg_field NumQSFPInterfaces;
	uvm_reg_field HSSI_CAPABILITY_num_channels;
	uvm_reg_field num_channels;
	uvm_reg_field HSSI_CAPABILITY_Num_channels_CSR_interface;
	uvm_reg_field Num_channels_CSR_interface;
	uvm_reg_field HSSI_CAPABILITY_Num_CSR_interface;
	uvm_reg_field Num_CSR_interface;
	rand uvm_reg_field HSSI_CTRL_Reserved;
	uvm_reg_field HSSI_STAT0_Chan3RxReady;
	uvm_reg_field Chan3RxReady;
	uvm_reg_field HSSI_STAT0_Chan3TxReady;
	uvm_reg_field Chan3TxReady;
	uvm_reg_field HSSI_STAT0_Chan3RxIsLockedToRef;
	uvm_reg_field Chan3RxIsLockedToRef;
	uvm_reg_field HSSI_STAT0_Chan3RxIsLockedToData;
	uvm_reg_field Chan3RxIsLockedToData;
	uvm_reg_field HSSI_STAT0_EChan3RxCalBusy;
	uvm_reg_field EChan3RxCalBusy;
	uvm_reg_field HSSI_STAT0_Chan3TxCalBusy;
	uvm_reg_field Chan3TxCalBusy;
	uvm_reg_field HSSI_STAT0_Chan3RxTransferReady;
	uvm_reg_field Chan3RxTransferReady;
	uvm_reg_field HSSI_STAT0_Chan3TxTransferReady;
	uvm_reg_field Chan3TxTransferReady;
	uvm_reg_field HSSI_STAT0_Chan3RxFifoReady;
	uvm_reg_field Chan3RxFifoReady;
	uvm_reg_field HSSI_STAT0_Chan3TxFifoReady;
	uvm_reg_field Chan3TxFifoReady;
	uvm_reg_field HSSI_STAT0_Chan3RxDigitalResetTimeout;
	uvm_reg_field Chan3RxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT0_Chan3TxDigitalResetTimeout;
	uvm_reg_field Chan3TxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT0_Chan3RxDigitalResetStat;
	uvm_reg_field Chan3RxDigitalResetStat;
	uvm_reg_field HSSI_STAT0_Chan3RxAnalogResetStat;
	uvm_reg_field Chan3RxAnalogResetStat;
	uvm_reg_field HSSI_STAT0_Chan3TxDigitalResetStat;
	uvm_reg_field Chan3TxDigitalResetStat;
	uvm_reg_field HSSI_STAT0_Chan3TxAnalogResetStat;
	uvm_reg_field Chan3TxAnalogResetStat;
	uvm_reg_field HSSI_STAT0_Chan2RxReady;
	uvm_reg_field Chan2RxReady;
	uvm_reg_field HSSI_STAT0_Chan2TxReady;
	uvm_reg_field Chan2TxReady;
	uvm_reg_field HSSI_STAT0_Chan2RxIsLockedToRef;
	uvm_reg_field Chan2RxIsLockedToRef;
	uvm_reg_field HSSI_STAT0_Chan2RxIsLockedToData;
	uvm_reg_field Chan2RxIsLockedToData;
	uvm_reg_field HSSI_STAT0_Chan2RxCalBusy;
	uvm_reg_field Chan2RxCalBusy;
	uvm_reg_field HSSI_STAT0_Chan2TxCalBusy;
	uvm_reg_field Chan2TxCalBusy;
	uvm_reg_field HSSI_STAT0_Chan2RxTransferReady;
	uvm_reg_field Chan2RxTransferReady;
	uvm_reg_field HSSI_STAT0_Chan2TxTransferReady;
	uvm_reg_field Chan2TxTransferReady;
	uvm_reg_field HSSI_STAT0_Chan2RxFifoReady;
	uvm_reg_field Chan2RxFifoReady;
	uvm_reg_field HSSI_STAT0_Chan2TxFifoReady;
	uvm_reg_field Chan2TxFifoReady;
	uvm_reg_field HSSI_STAT0_Chan2RxDigitalResetTimeout;
	uvm_reg_field Chan2RxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT0_Chan2TxDigitalResetTimeout;
	uvm_reg_field Chan2TxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT0_Chan2RxDigitalResetStat;
	uvm_reg_field Chan2RxDigitalResetStat;
	uvm_reg_field HSSI_STAT0_Chan2RxAnalogResetStat;
	uvm_reg_field Chan2RxAnalogResetStat;
	uvm_reg_field HSSI_STAT0_Chan2TxDigitalResetStat;
	uvm_reg_field Chan2TxDigitalResetStat;
	uvm_reg_field HSSI_STAT0_Chan2TxAnalogResetStat;
	uvm_reg_field Chan2TxAnalogResetStat;
	uvm_reg_field HSSI_STAT0_Chan1RxReady;
	uvm_reg_field Chan1RxReady;
	uvm_reg_field HSSI_STAT0_Chan1TxReady;
	uvm_reg_field Chan1TxReady;
	uvm_reg_field HSSI_STAT0_Chan1RxIsLockedToRef;
	uvm_reg_field Chan1RxIsLockedToRef;
	uvm_reg_field HSSI_STAT0_Chan1RxIsLockedToData;
	uvm_reg_field Chan1RxIsLockedToData;
	uvm_reg_field HSSI_STAT0_Chan1RxCalBusy;
	uvm_reg_field Chan1RxCalBusy;
	uvm_reg_field HSSI_STAT0_Chan1TxCalBusy;
	uvm_reg_field HSSI_STAT0_Chan1RxTransferReady;
	uvm_reg_field Chan1RxTransferReady;
	uvm_reg_field HSSI_STAT0_Chan1TxTransferReady;
	uvm_reg_field Chan1TxTransferReady;
	uvm_reg_field HSSI_STAT0_Chan1RxFifoReady;
	uvm_reg_field Chan1RxFifoReady;
	uvm_reg_field HSSI_STAT0_Chan1TxFifoReady;
	uvm_reg_field Chan1TxFifoReady;
	uvm_reg_field HSSI_STAT0_Chan1RxDigitalResetTimeout;
	uvm_reg_field Chan1RxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT0_Chan1TxDigitalResetTimeout;
	uvm_reg_field Chan1TxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT0_Chan1RxDigitalResetStat;
	uvm_reg_field Chan1RxDigitalResetStat;
	uvm_reg_field HSSI_STAT0_Chan1RxAnalogResetStat;
	uvm_reg_field Chan1RxAnalogResetStat;
	uvm_reg_field HSSI_STAT0_Chan1TxDigitalResetStat;
	uvm_reg_field Chan1TxDigitalResetStat;
	uvm_reg_field HSSI_STAT0_Chan1TxAnalogResetStat;
	uvm_reg_field Chan1TxAnalogResetStat;
	uvm_reg_field HSSI_STAT0_Chan0RxReady;
	uvm_reg_field Chan0RxReady;
	uvm_reg_field HSSI_STAT0_Chan0TxReady;
	uvm_reg_field Chan0TxReady;
	uvm_reg_field HSSI_STAT0_Chan0RxIsLockedToRef;
	uvm_reg_field Chan0RxIsLockedToRef;
	uvm_reg_field HSSI_STAT0_Chan0RxIsLockedToData;
	uvm_reg_field Chan0RxIsLockedToData;
	uvm_reg_field HSSI_STAT0_Chan0RxCalBusy;
	uvm_reg_field Chan0RxCalBusy;
	uvm_reg_field HSSI_STAT0_Chan0TxCalBusy;
	uvm_reg_field Chan0TxCalBusy;
	uvm_reg_field HSSI_STAT0_Chan0RxTransferReady;
	uvm_reg_field Chan0RxTransferReady;
	uvm_reg_field HSSI_STAT0_Chan0TxTransferReady;
	uvm_reg_field Chan0TxTransferReady;
	uvm_reg_field HSSI_STAT0_Chan0RxFifoReady;
	uvm_reg_field Chan0RxFifoReady;
	uvm_reg_field HSSI_STAT0_Chan0TxFifoReady;
	uvm_reg_field Chan0TxFifoReady;
	uvm_reg_field HSSI_STAT0_Chan0RxDigitalResetTimeout;
	uvm_reg_field Chan0RxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT0_Chan0TxDigitalResetTimeout;
	uvm_reg_field Chan0TxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT0_Chan0RxDigitalResetStat;
	uvm_reg_field Chan0RxDigitalResetStat;
	uvm_reg_field HSSI_STAT0_Chan0RxAnalogResetStat;
	uvm_reg_field Chan0RxAnalogResetStat;
	uvm_reg_field HSSI_STAT0_Chan0TxDigitalResetStat;
	uvm_reg_field Chan0TxDigitalResetStat;
	uvm_reg_field HSSI_STAT0_Chan0TxAnalogResetStat;
	uvm_reg_field Chan0TxAnalogResetStat;
	uvm_reg_field HSSI_STAT1_Chan7RxReady;
	uvm_reg_field Chan7RxReady;
	uvm_reg_field HSSI_STAT1_Chan7TxReady;
	uvm_reg_field Chan7TxReady;
	uvm_reg_field HSSI_STAT1_Chan7RxIsLockedToRef;
	uvm_reg_field Chan7RxIsLockedToRef;
	uvm_reg_field HSSI_STAT1_Chan7RxIsLockedToData;
	uvm_reg_field Chan7RxIsLockedToData;
	uvm_reg_field HSSI_STAT1_EChan7RxCalBusy;
	uvm_reg_field EChan7RxCalBusy;
	uvm_reg_field HSSI_STAT1_Chan7TxCalBusy;
	uvm_reg_field Chan7TxCalBusy;
	uvm_reg_field HSSI_STAT1_Chan7RxTransferReady;
	uvm_reg_field Chan7RxTransferReady;
	uvm_reg_field HSSI_STAT1_Chan7TxTransferReady;
	uvm_reg_field Chan7TxTransferReady;
	uvm_reg_field HSSI_STAT1_Chan7RxFifoReady;
	uvm_reg_field Chan7RxFifoReady;
	uvm_reg_field HSSI_STAT1_Chan7TxFifoReady;
	uvm_reg_field Chan7TxFifoReady;
	uvm_reg_field HSSI_STAT1_Chan7RxDigitalResetTimeout;
	uvm_reg_field Chan7RxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT1_Chan7TxDigitalResetTimeout;
	uvm_reg_field Chan7TxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT1_Chan7RxDigitalResetStat;
	uvm_reg_field Chan7RxDigitalResetStat;
	uvm_reg_field HSSI_STAT1_Chan7RxAnalogResetStat;
	uvm_reg_field Chan7RxAnalogResetStat;
	uvm_reg_field HSSI_STAT1_Chan7TxDigitalResetStat;
	uvm_reg_field Chan7TxDigitalResetStat;
	uvm_reg_field HSSI_STAT1_Chan7TxAnalogResetStat;
	uvm_reg_field Chan7TxAnalogResetStat;
	uvm_reg_field HSSI_STAT1_Chan6RxReady;
	uvm_reg_field Chan6RxReady;
	uvm_reg_field HSSI_STAT1_Chan6TxReady;
	uvm_reg_field Chan6TxReady;
	uvm_reg_field HSSI_STAT1_Chan6RxIsLockedToRef;
	uvm_reg_field Chan6RxIsLockedToRef;
	uvm_reg_field HSSI_STAT1_Chan6RxIsLockedToData;
	uvm_reg_field Chan6RxIsLockedToData;
	uvm_reg_field HSSI_STAT1_Chan6RxCalBusy;
	uvm_reg_field Chan6RxCalBusy;
	uvm_reg_field HSSI_STAT1_Chan6TxCalBusy;
	uvm_reg_field Chan6TxCalBusy;
	uvm_reg_field HSSI_STAT1_Chan6RxTransferReady;
	uvm_reg_field Chan6RxTransferReady;
	uvm_reg_field HSSI_STAT1_Chan6TxTransferReady;
	uvm_reg_field Chan6TxTransferReady;
	uvm_reg_field HSSI_STAT1_Chan6RxFifoReady;
	uvm_reg_field Chan6RxFifoReady;
	uvm_reg_field HSSI_STAT1_Chan6TxFifoReady;
	uvm_reg_field Chan6TxFifoReady;
	uvm_reg_field HSSI_STAT1_Chan6RxDigitalResetTimeout;
	uvm_reg_field Chan6RxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT1_Chan6TxDigitalResetTimeout;
	uvm_reg_field Chan6TxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT1_Chan6RxDigitalResetStat;
	uvm_reg_field Chan6RxDigitalResetStat;
	uvm_reg_field HSSI_STAT1_Chan6RxAnalogResetStat;
	uvm_reg_field Chan6RxAnalogResetStat;
	uvm_reg_field HSSI_STAT1_Chan6TxDigitalResetStat;
	uvm_reg_field Chan6TxDigitalResetStat;
	uvm_reg_field HSSI_STAT1_Chan6TxAnalogResetStat;
	uvm_reg_field Chan6TxAnalogResetStat;
	uvm_reg_field HSSI_STAT1_Chan5RxReady;
	uvm_reg_field Chan5RxReady;
	uvm_reg_field HSSI_STAT1_Chan5TxReady;
	uvm_reg_field Chan5TxReady;
	uvm_reg_field HSSI_STAT1_Chan5RxIsLockedToRef;
	uvm_reg_field Chan5RxIsLockedToRef;
	uvm_reg_field HSSI_STAT1_Chan5RxIsLockedToData;
	uvm_reg_field Chan5RxIsLockedToData;
	uvm_reg_field HSSI_STAT1_Chan5RxCalBusy;
	uvm_reg_field Chan5RxCalBusy;
	uvm_reg_field HSSI_STAT1_Chan1TxCalBusy;
	uvm_reg_field HSSI_STAT1_Chan5RxTransferReady;
	uvm_reg_field Chan5RxTransferReady;
	uvm_reg_field HSSI_STAT1_Chan5TxTransferReady;
	uvm_reg_field Chan5TxTransferReady;
	uvm_reg_field HSSI_STAT1_Chan5RxFifoReady;
	uvm_reg_field Chan5RxFifoReady;
	uvm_reg_field HSSI_STAT1_Chan5TxFifoReady;
	uvm_reg_field Chan5TxFifoReady;
	uvm_reg_field HSSI_STAT1_Chan5RxDigitalResetTimeout;
	uvm_reg_field Chan5RxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT1_Chan5TxDigitalResetTimeout;
	uvm_reg_field Chan5TxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT1_Chan5RxDigitalResetStat;
	uvm_reg_field Chan5RxDigitalResetStat;
	uvm_reg_field HSSI_STAT1_Chan5RxAnalogResetStat;
	uvm_reg_field Chan5RxAnalogResetStat;
	uvm_reg_field HSSI_STAT1_Chan5TxDigitalResetStat;
	uvm_reg_field Chan5TxDigitalResetStat;
	uvm_reg_field HSSI_STAT1_Chan5TxAnalogResetStat;
	uvm_reg_field Chan5TxAnalogResetStat;
	uvm_reg_field HSSI_STAT1_Chan4RxReady;
	uvm_reg_field Chan4RxReady;
	uvm_reg_field HSSI_STAT1_Chan4TxReady;
	uvm_reg_field Chan4TxReady;
	uvm_reg_field HSSI_STAT1_Chan4RxIsLockedToRef;
	uvm_reg_field Chan4RxIsLockedToRef;
	uvm_reg_field HSSI_STAT1_Chan4RxIsLockedToData;
	uvm_reg_field Chan4RxIsLockedToData;
	uvm_reg_field HSSI_STAT1_Chan4RxCalBusy;
	uvm_reg_field Chan4RxCalBusy;
	uvm_reg_field HSSI_STAT1_Chan4TxCalBusy;
	uvm_reg_field Chan4TxCalBusy;
	uvm_reg_field HSSI_STAT1_Chan4RxTransferReady;
	uvm_reg_field Chan4RxTransferReady;
	uvm_reg_field HSSI_STAT1_Chan4TxTransferReady;
	uvm_reg_field Chan4TxTransferReady;
	uvm_reg_field HSSI_STAT1_Chan4RxFifoReady;
	uvm_reg_field Chan4RxFifoReady;
	uvm_reg_field HSSI_STAT1_Chan4TxFifoReady;
	uvm_reg_field Chan4TxFifoReady;
	uvm_reg_field HSSI_STAT1_Chan4RxDigitalResetTimeout;
	uvm_reg_field Chan4RxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT1_Chan4TxDigitalResetTimeout;
	uvm_reg_field Chan4TxDigitalResetTimeout;
	uvm_reg_field HSSI_STAT1_Chan4RxDigitalResetStat;
	uvm_reg_field Chan4RxDigitalResetStat;
	uvm_reg_field HSSI_STAT1_Chan4RxAnalogResetStat;
	uvm_reg_field Chan4RxAnalogResetStat;
	uvm_reg_field HSSI_STAT1_Chan4TxDigitalResetStat;
	uvm_reg_field Chan4TxDigitalResetStat;
	uvm_reg_field HSSI_STAT1_Chan4TxAnalogResetStat;
	uvm_reg_field Chan4TxAnalogResetStat;
	rand uvm_reg_field HSSI_RCFG_CMD0_Reserved;
	rand uvm_reg_field HSSI_RCFG_CMD0_XcvrRcfgAddr;
	rand uvm_reg_field XcvrRcfgAddr;
	rand uvm_reg_field HSSI_RCFG_CMD0_Reserved_1;
	rand uvm_reg_field Reserved_1;
	uvm_reg_field HSSI_RCFG_CMD0_XcvrRcfgAck;
	uvm_reg_field XcvrRcfgAck;
	rand uvm_reg_field HSSI_RCFG_CMD0_XcvrRcfgCmdStatus;
	rand uvm_reg_field XcvrRcfgCmdStatus;
	rand uvm_reg_field HSSI_RCFG_DATA0_XcvrRcfgWrData;
	rand uvm_reg_field XcvrRcfgWrData;
	uvm_reg_field HSSI_RCFG_DATA0_XcvrRcfgRdData;
	uvm_reg_field XcvrRcfgRdData;
	rand uvm_reg_field HSSI_SCRATCHPAD_Scrathpad;
	rand uvm_reg_field Scrathpad;

	function new(string name = "hssi_ss_csr");
		super.new(name, build_coverage(UVM_NO_COVERAGE));
	endfunction: new

   virtual function void build();
      this.default_map = create_map("", 0, 8, UVM_LITTLE_ENDIAN, 0);
      this.HSSI_DFH = ral_reg_hssi_ss_csr_HSSI_DFH::type_id::create("HSSI_DFH",,get_full_name());
      this.HSSI_DFH.configure(this, null, "");
      this.HSSI_DFH.build();
      this.default_map.add_reg(this.HSSI_DFH, `UVM_REG_ADDR_WIDTH'h0, "RW", 0);
		this.HSSI_DFH_FeatureType = this.HSSI_DFH.FeatureType;
		this.FeatureType = this.HSSI_DFH.FeatureType;
		this.HSSI_DFH_Reserved = this.HSSI_DFH.Reserved;
		this.HSSI_DFH_EOL = this.HSSI_DFH.EOL;
		this.EOL = this.HSSI_DFH.EOL;
		this.HSSI_DFH_NextDfhByteOffset = this.HSSI_DFH.NextDfhByteOffset;
		this.NextDfhByteOffset = this.HSSI_DFH.NextDfhByteOffset;
		this.HSSI_DFH_FeatureRevision = this.HSSI_DFH.FeatureRevision;
		this.FeatureRevision = this.HSSI_DFH.FeatureRevision;
		this.HSSI_DFH_FeatureId = this.HSSI_DFH.FeatureId;
		this.FeatureId = this.HSSI_DFH.FeatureId;
      this.HSSI_CAPABILITY = ral_reg_hssi_ss_csr_HSSI_CAPABILITY::type_id::create("HSSI_CAPABILITY",,get_full_name());
      this.HSSI_CAPABILITY.configure(this, null, "");
      this.HSSI_CAPABILITY.build();
      this.default_map.add_reg(this.HSSI_CAPABILITY, `UVM_REG_ADDR_WIDTH'h8, "RW", 0);
		this.HSSI_CAPABILITY_Reserved = this.HSSI_CAPABILITY.Reserved;
		this.HSSI_CAPABILITY_NumQSFPInterfaces = this.HSSI_CAPABILITY.NumQSFPInterfaces;
		this.NumQSFPInterfaces = this.HSSI_CAPABILITY.NumQSFPInterfaces;
		this.HSSI_CAPABILITY_num_channels = this.HSSI_CAPABILITY.num_channels;
		this.num_channels = this.HSSI_CAPABILITY.num_channels;
		this.HSSI_CAPABILITY_Num_channels_CSR_interface = this.HSSI_CAPABILITY.Num_channels_CSR_interface;
		this.Num_channels_CSR_interface = this.HSSI_CAPABILITY.Num_channels_CSR_interface;
		this.HSSI_CAPABILITY_Num_CSR_interface = this.HSSI_CAPABILITY.Num_CSR_interface;
		this.Num_CSR_interface = this.HSSI_CAPABILITY.Num_CSR_interface;
      this.HSSI_CTRL = ral_reg_hssi_ss_csr_HSSI_CTRL::type_id::create("HSSI_CTRL",,get_full_name());
      this.HSSI_CTRL.configure(this, null, "");
      this.HSSI_CTRL.build();
      this.default_map.add_reg(this.HSSI_CTRL, `UVM_REG_ADDR_WIDTH'h10, "RW", 0);
		this.HSSI_CTRL_Reserved = this.HSSI_CTRL.Reserved;
      this.HSSI_STAT0 = ral_reg_hssi_ss_csr_HSSI_STAT0::type_id::create("HSSI_STAT0",,get_full_name());
      this.HSSI_STAT0.configure(this, null, "");
      this.HSSI_STAT0.build();
      this.default_map.add_reg(this.HSSI_STAT0, `UVM_REG_ADDR_WIDTH'h18, "RO", 0);
		this.HSSI_STAT0_Chan3RxReady = this.HSSI_STAT0.Chan3RxReady;
		this.Chan3RxReady = this.HSSI_STAT0.Chan3RxReady;
		this.HSSI_STAT0_Chan3TxReady = this.HSSI_STAT0.Chan3TxReady;
		this.Chan3TxReady = this.HSSI_STAT0.Chan3TxReady;
		this.HSSI_STAT0_Chan3RxIsLockedToRef = this.HSSI_STAT0.Chan3RxIsLockedToRef;
		this.Chan3RxIsLockedToRef = this.HSSI_STAT0.Chan3RxIsLockedToRef;
		this.HSSI_STAT0_Chan3RxIsLockedToData = this.HSSI_STAT0.Chan3RxIsLockedToData;
		this.Chan3RxIsLockedToData = this.HSSI_STAT0.Chan3RxIsLockedToData;
		this.HSSI_STAT0_EChan3RxCalBusy = this.HSSI_STAT0.EChan3RxCalBusy;
		this.EChan3RxCalBusy = this.HSSI_STAT0.EChan3RxCalBusy;
		this.HSSI_STAT0_Chan3TxCalBusy = this.HSSI_STAT0.Chan3TxCalBusy;
		this.Chan3TxCalBusy = this.HSSI_STAT0.Chan3TxCalBusy;
		this.HSSI_STAT0_Chan3RxTransferReady = this.HSSI_STAT0.Chan3RxTransferReady;
		this.Chan3RxTransferReady = this.HSSI_STAT0.Chan3RxTransferReady;
		this.HSSI_STAT0_Chan3TxTransferReady = this.HSSI_STAT0.Chan3TxTransferReady;
		this.Chan3TxTransferReady = this.HSSI_STAT0.Chan3TxTransferReady;
		this.HSSI_STAT0_Chan3RxFifoReady = this.HSSI_STAT0.Chan3RxFifoReady;
		this.Chan3RxFifoReady = this.HSSI_STAT0.Chan3RxFifoReady;
		this.HSSI_STAT0_Chan3TxFifoReady = this.HSSI_STAT0.Chan3TxFifoReady;
		this.Chan3TxFifoReady = this.HSSI_STAT0.Chan3TxFifoReady;
		this.HSSI_STAT0_Chan3RxDigitalResetTimeout = this.HSSI_STAT0.Chan3RxDigitalResetTimeout;
		this.Chan3RxDigitalResetTimeout = this.HSSI_STAT0.Chan3RxDigitalResetTimeout;
		this.HSSI_STAT0_Chan3TxDigitalResetTimeout = this.HSSI_STAT0.Chan3TxDigitalResetTimeout;
		this.Chan3TxDigitalResetTimeout = this.HSSI_STAT0.Chan3TxDigitalResetTimeout;
		this.HSSI_STAT0_Chan3RxDigitalResetStat = this.HSSI_STAT0.Chan3RxDigitalResetStat;
		this.Chan3RxDigitalResetStat = this.HSSI_STAT0.Chan3RxDigitalResetStat;
		this.HSSI_STAT0_Chan3RxAnalogResetStat = this.HSSI_STAT0.Chan3RxAnalogResetStat;
		this.Chan3RxAnalogResetStat = this.HSSI_STAT0.Chan3RxAnalogResetStat;
		this.HSSI_STAT0_Chan3TxDigitalResetStat = this.HSSI_STAT0.Chan3TxDigitalResetStat;
		this.Chan3TxDigitalResetStat = this.HSSI_STAT0.Chan3TxDigitalResetStat;
		this.HSSI_STAT0_Chan3TxAnalogResetStat = this.HSSI_STAT0.Chan3TxAnalogResetStat;
		this.Chan3TxAnalogResetStat = this.HSSI_STAT0.Chan3TxAnalogResetStat;
		this.HSSI_STAT0_Chan2RxReady = this.HSSI_STAT0.Chan2RxReady;
		this.Chan2RxReady = this.HSSI_STAT0.Chan2RxReady;
		this.HSSI_STAT0_Chan2TxReady = this.HSSI_STAT0.Chan2TxReady;
		this.Chan2TxReady = this.HSSI_STAT0.Chan2TxReady;
		this.HSSI_STAT0_Chan2RxIsLockedToRef = this.HSSI_STAT0.Chan2RxIsLockedToRef;
		this.Chan2RxIsLockedToRef = this.HSSI_STAT0.Chan2RxIsLockedToRef;
		this.HSSI_STAT0_Chan2RxIsLockedToData = this.HSSI_STAT0.Chan2RxIsLockedToData;
		this.Chan2RxIsLockedToData = this.HSSI_STAT0.Chan2RxIsLockedToData;
		this.HSSI_STAT0_Chan2RxCalBusy = this.HSSI_STAT0.Chan2RxCalBusy;
		this.Chan2RxCalBusy = this.HSSI_STAT0.Chan2RxCalBusy;
		this.HSSI_STAT0_Chan2TxCalBusy = this.HSSI_STAT0.Chan2TxCalBusy;
		this.Chan2TxCalBusy = this.HSSI_STAT0.Chan2TxCalBusy;
		this.HSSI_STAT0_Chan2RxTransferReady = this.HSSI_STAT0.Chan2RxTransferReady;
		this.Chan2RxTransferReady = this.HSSI_STAT0.Chan2RxTransferReady;
		this.HSSI_STAT0_Chan2TxTransferReady = this.HSSI_STAT0.Chan2TxTransferReady;
		this.Chan2TxTransferReady = this.HSSI_STAT0.Chan2TxTransferReady;
		this.HSSI_STAT0_Chan2RxFifoReady = this.HSSI_STAT0.Chan2RxFifoReady;
		this.Chan2RxFifoReady = this.HSSI_STAT0.Chan2RxFifoReady;
		this.HSSI_STAT0_Chan2TxFifoReady = this.HSSI_STAT0.Chan2TxFifoReady;
		this.Chan2TxFifoReady = this.HSSI_STAT0.Chan2TxFifoReady;
		this.HSSI_STAT0_Chan2RxDigitalResetTimeout = this.HSSI_STAT0.Chan2RxDigitalResetTimeout;
		this.Chan2RxDigitalResetTimeout = this.HSSI_STAT0.Chan2RxDigitalResetTimeout;
		this.HSSI_STAT0_Chan2TxDigitalResetTimeout = this.HSSI_STAT0.Chan2TxDigitalResetTimeout;
		this.Chan2TxDigitalResetTimeout = this.HSSI_STAT0.Chan2TxDigitalResetTimeout;
		this.HSSI_STAT0_Chan2RxDigitalResetStat = this.HSSI_STAT0.Chan2RxDigitalResetStat;
		this.Chan2RxDigitalResetStat = this.HSSI_STAT0.Chan2RxDigitalResetStat;
		this.HSSI_STAT0_Chan2RxAnalogResetStat = this.HSSI_STAT0.Chan2RxAnalogResetStat;
		this.Chan2RxAnalogResetStat = this.HSSI_STAT0.Chan2RxAnalogResetStat;
		this.HSSI_STAT0_Chan2TxDigitalResetStat = this.HSSI_STAT0.Chan2TxDigitalResetStat;
		this.Chan2TxDigitalResetStat = this.HSSI_STAT0.Chan2TxDigitalResetStat;
		this.HSSI_STAT0_Chan2TxAnalogResetStat = this.HSSI_STAT0.Chan2TxAnalogResetStat;
		this.Chan2TxAnalogResetStat = this.HSSI_STAT0.Chan2TxAnalogResetStat;
		this.HSSI_STAT0_Chan1RxReady = this.HSSI_STAT0.Chan1RxReady;
		this.Chan1RxReady = this.HSSI_STAT0.Chan1RxReady;
		this.HSSI_STAT0_Chan1TxReady = this.HSSI_STAT0.Chan1TxReady;
		this.Chan1TxReady = this.HSSI_STAT0.Chan1TxReady;
		this.HSSI_STAT0_Chan1RxIsLockedToRef = this.HSSI_STAT0.Chan1RxIsLockedToRef;
		this.Chan1RxIsLockedToRef = this.HSSI_STAT0.Chan1RxIsLockedToRef;
		this.HSSI_STAT0_Chan1RxIsLockedToData = this.HSSI_STAT0.Chan1RxIsLockedToData;
		this.Chan1RxIsLockedToData = this.HSSI_STAT0.Chan1RxIsLockedToData;
		this.HSSI_STAT0_Chan1RxCalBusy = this.HSSI_STAT0.Chan1RxCalBusy;
		this.Chan1RxCalBusy = this.HSSI_STAT0.Chan1RxCalBusy;
		this.HSSI_STAT0_Chan1TxCalBusy = this.HSSI_STAT0.Chan1TxCalBusy;
		this.HSSI_STAT0_Chan1RxTransferReady = this.HSSI_STAT0.Chan1RxTransferReady;
		this.Chan1RxTransferReady = this.HSSI_STAT0.Chan1RxTransferReady;
		this.HSSI_STAT0_Chan1TxTransferReady = this.HSSI_STAT0.Chan1TxTransferReady;
		this.Chan1TxTransferReady = this.HSSI_STAT0.Chan1TxTransferReady;
		this.HSSI_STAT0_Chan1RxFifoReady = this.HSSI_STAT0.Chan1RxFifoReady;
		this.Chan1RxFifoReady = this.HSSI_STAT0.Chan1RxFifoReady;
		this.HSSI_STAT0_Chan1TxFifoReady = this.HSSI_STAT0.Chan1TxFifoReady;
		this.Chan1TxFifoReady = this.HSSI_STAT0.Chan1TxFifoReady;
		this.HSSI_STAT0_Chan1RxDigitalResetTimeout = this.HSSI_STAT0.Chan1RxDigitalResetTimeout;
		this.Chan1RxDigitalResetTimeout = this.HSSI_STAT0.Chan1RxDigitalResetTimeout;
		this.HSSI_STAT0_Chan1TxDigitalResetTimeout = this.HSSI_STAT0.Chan1TxDigitalResetTimeout;
		this.Chan1TxDigitalResetTimeout = this.HSSI_STAT0.Chan1TxDigitalResetTimeout;
		this.HSSI_STAT0_Chan1RxDigitalResetStat = this.HSSI_STAT0.Chan1RxDigitalResetStat;
		this.Chan1RxDigitalResetStat = this.HSSI_STAT0.Chan1RxDigitalResetStat;
		this.HSSI_STAT0_Chan1RxAnalogResetStat = this.HSSI_STAT0.Chan1RxAnalogResetStat;
		this.Chan1RxAnalogResetStat = this.HSSI_STAT0.Chan1RxAnalogResetStat;
		this.HSSI_STAT0_Chan1TxDigitalResetStat = this.HSSI_STAT0.Chan1TxDigitalResetStat;
		this.Chan1TxDigitalResetStat = this.HSSI_STAT0.Chan1TxDigitalResetStat;
		this.HSSI_STAT0_Chan1TxAnalogResetStat = this.HSSI_STAT0.Chan1TxAnalogResetStat;
		this.Chan1TxAnalogResetStat = this.HSSI_STAT0.Chan1TxAnalogResetStat;
		this.HSSI_STAT0_Chan0RxReady = this.HSSI_STAT0.Chan0RxReady;
		this.Chan0RxReady = this.HSSI_STAT0.Chan0RxReady;
		this.HSSI_STAT0_Chan0TxReady = this.HSSI_STAT0.Chan0TxReady;
		this.Chan0TxReady = this.HSSI_STAT0.Chan0TxReady;
		this.HSSI_STAT0_Chan0RxIsLockedToRef = this.HSSI_STAT0.Chan0RxIsLockedToRef;
		this.Chan0RxIsLockedToRef = this.HSSI_STAT0.Chan0RxIsLockedToRef;
		this.HSSI_STAT0_Chan0RxIsLockedToData = this.HSSI_STAT0.Chan0RxIsLockedToData;
		this.Chan0RxIsLockedToData = this.HSSI_STAT0.Chan0RxIsLockedToData;
		this.HSSI_STAT0_Chan0RxCalBusy = this.HSSI_STAT0.Chan0RxCalBusy;
		this.Chan0RxCalBusy = this.HSSI_STAT0.Chan0RxCalBusy;
		this.HSSI_STAT0_Chan0TxCalBusy = this.HSSI_STAT0.Chan0TxCalBusy;
		this.Chan0TxCalBusy = this.HSSI_STAT0.Chan0TxCalBusy;
		this.HSSI_STAT0_Chan0RxTransferReady = this.HSSI_STAT0.Chan0RxTransferReady;
		this.Chan0RxTransferReady = this.HSSI_STAT0.Chan0RxTransferReady;
		this.HSSI_STAT0_Chan0TxTransferReady = this.HSSI_STAT0.Chan0TxTransferReady;
		this.Chan0TxTransferReady = this.HSSI_STAT0.Chan0TxTransferReady;
		this.HSSI_STAT0_Chan0RxFifoReady = this.HSSI_STAT0.Chan0RxFifoReady;
		this.Chan0RxFifoReady = this.HSSI_STAT0.Chan0RxFifoReady;
		this.HSSI_STAT0_Chan0TxFifoReady = this.HSSI_STAT0.Chan0TxFifoReady;
		this.Chan0TxFifoReady = this.HSSI_STAT0.Chan0TxFifoReady;
		this.HSSI_STAT0_Chan0RxDigitalResetTimeout = this.HSSI_STAT0.Chan0RxDigitalResetTimeout;
		this.Chan0RxDigitalResetTimeout = this.HSSI_STAT0.Chan0RxDigitalResetTimeout;
		this.HSSI_STAT0_Chan0TxDigitalResetTimeout = this.HSSI_STAT0.Chan0TxDigitalResetTimeout;
		this.Chan0TxDigitalResetTimeout = this.HSSI_STAT0.Chan0TxDigitalResetTimeout;
		this.HSSI_STAT0_Chan0RxDigitalResetStat = this.HSSI_STAT0.Chan0RxDigitalResetStat;
		this.Chan0RxDigitalResetStat = this.HSSI_STAT0.Chan0RxDigitalResetStat;
		this.HSSI_STAT0_Chan0RxAnalogResetStat = this.HSSI_STAT0.Chan0RxAnalogResetStat;
		this.Chan0RxAnalogResetStat = this.HSSI_STAT0.Chan0RxAnalogResetStat;
		this.HSSI_STAT0_Chan0TxDigitalResetStat = this.HSSI_STAT0.Chan0TxDigitalResetStat;
		this.Chan0TxDigitalResetStat = this.HSSI_STAT0.Chan0TxDigitalResetStat;
		this.HSSI_STAT0_Chan0TxAnalogResetStat = this.HSSI_STAT0.Chan0TxAnalogResetStat;
		this.Chan0TxAnalogResetStat = this.HSSI_STAT0.Chan0TxAnalogResetStat;
      this.HSSI_STAT1 = ral_reg_hssi_ss_csr_HSSI_STAT1::type_id::create("HSSI_STAT1",,get_full_name());
      this.HSSI_STAT1.configure(this, null, "");
      this.HSSI_STAT1.build();
      this.default_map.add_reg(this.HSSI_STAT1, `UVM_REG_ADDR_WIDTH'h20, "RO", 0);
		this.HSSI_STAT1_Chan7RxReady = this.HSSI_STAT1.Chan7RxReady;
		this.Chan7RxReady = this.HSSI_STAT1.Chan7RxReady;
		this.HSSI_STAT1_Chan7TxReady = this.HSSI_STAT1.Chan7TxReady;
		this.Chan7TxReady = this.HSSI_STAT1.Chan7TxReady;
		this.HSSI_STAT1_Chan7RxIsLockedToRef = this.HSSI_STAT1.Chan7RxIsLockedToRef;
		this.Chan7RxIsLockedToRef = this.HSSI_STAT1.Chan7RxIsLockedToRef;
		this.HSSI_STAT1_Chan7RxIsLockedToData = this.HSSI_STAT1.Chan7RxIsLockedToData;
		this.Chan7RxIsLockedToData = this.HSSI_STAT1.Chan7RxIsLockedToData;
		this.HSSI_STAT1_EChan7RxCalBusy = this.HSSI_STAT1.EChan7RxCalBusy;
		this.EChan7RxCalBusy = this.HSSI_STAT1.EChan7RxCalBusy;
		this.HSSI_STAT1_Chan7TxCalBusy = this.HSSI_STAT1.Chan7TxCalBusy;
		this.Chan7TxCalBusy = this.HSSI_STAT1.Chan7TxCalBusy;
		this.HSSI_STAT1_Chan7RxTransferReady = this.HSSI_STAT1.Chan7RxTransferReady;
		this.Chan7RxTransferReady = this.HSSI_STAT1.Chan7RxTransferReady;
		this.HSSI_STAT1_Chan7TxTransferReady = this.HSSI_STAT1.Chan7TxTransferReady;
		this.Chan7TxTransferReady = this.HSSI_STAT1.Chan7TxTransferReady;
		this.HSSI_STAT1_Chan7RxFifoReady = this.HSSI_STAT1.Chan7RxFifoReady;
		this.Chan7RxFifoReady = this.HSSI_STAT1.Chan7RxFifoReady;
		this.HSSI_STAT1_Chan7TxFifoReady = this.HSSI_STAT1.Chan7TxFifoReady;
		this.Chan7TxFifoReady = this.HSSI_STAT1.Chan7TxFifoReady;
		this.HSSI_STAT1_Chan7RxDigitalResetTimeout = this.HSSI_STAT1.Chan7RxDigitalResetTimeout;
		this.Chan7RxDigitalResetTimeout = this.HSSI_STAT1.Chan7RxDigitalResetTimeout;
		this.HSSI_STAT1_Chan7TxDigitalResetTimeout = this.HSSI_STAT1.Chan7TxDigitalResetTimeout;
		this.Chan7TxDigitalResetTimeout = this.HSSI_STAT1.Chan7TxDigitalResetTimeout;
		this.HSSI_STAT1_Chan7RxDigitalResetStat = this.HSSI_STAT1.Chan7RxDigitalResetStat;
		this.Chan7RxDigitalResetStat = this.HSSI_STAT1.Chan7RxDigitalResetStat;
		this.HSSI_STAT1_Chan7RxAnalogResetStat = this.HSSI_STAT1.Chan7RxAnalogResetStat;
		this.Chan7RxAnalogResetStat = this.HSSI_STAT1.Chan7RxAnalogResetStat;
		this.HSSI_STAT1_Chan7TxDigitalResetStat = this.HSSI_STAT1.Chan7TxDigitalResetStat;
		this.Chan7TxDigitalResetStat = this.HSSI_STAT1.Chan7TxDigitalResetStat;
		this.HSSI_STAT1_Chan7TxAnalogResetStat = this.HSSI_STAT1.Chan7TxAnalogResetStat;
		this.Chan7TxAnalogResetStat = this.HSSI_STAT1.Chan7TxAnalogResetStat;
		this.HSSI_STAT1_Chan6RxReady = this.HSSI_STAT1.Chan6RxReady;
		this.Chan6RxReady = this.HSSI_STAT1.Chan6RxReady;
		this.HSSI_STAT1_Chan6TxReady = this.HSSI_STAT1.Chan6TxReady;
		this.Chan6TxReady = this.HSSI_STAT1.Chan6TxReady;
		this.HSSI_STAT1_Chan6RxIsLockedToRef = this.HSSI_STAT1.Chan6RxIsLockedToRef;
		this.Chan6RxIsLockedToRef = this.HSSI_STAT1.Chan6RxIsLockedToRef;
		this.HSSI_STAT1_Chan6RxIsLockedToData = this.HSSI_STAT1.Chan6RxIsLockedToData;
		this.Chan6RxIsLockedToData = this.HSSI_STAT1.Chan6RxIsLockedToData;
		this.HSSI_STAT1_Chan6RxCalBusy = this.HSSI_STAT1.Chan6RxCalBusy;
		this.Chan6RxCalBusy = this.HSSI_STAT1.Chan6RxCalBusy;
		this.HSSI_STAT1_Chan6TxCalBusy = this.HSSI_STAT1.Chan6TxCalBusy;
		this.Chan6TxCalBusy = this.HSSI_STAT1.Chan6TxCalBusy;
		this.HSSI_STAT1_Chan6RxTransferReady = this.HSSI_STAT1.Chan6RxTransferReady;
		this.Chan6RxTransferReady = this.HSSI_STAT1.Chan6RxTransferReady;
		this.HSSI_STAT1_Chan6TxTransferReady = this.HSSI_STAT1.Chan6TxTransferReady;
		this.Chan6TxTransferReady = this.HSSI_STAT1.Chan6TxTransferReady;
		this.HSSI_STAT1_Chan6RxFifoReady = this.HSSI_STAT1.Chan6RxFifoReady;
		this.Chan6RxFifoReady = this.HSSI_STAT1.Chan6RxFifoReady;
		this.HSSI_STAT1_Chan6TxFifoReady = this.HSSI_STAT1.Chan6TxFifoReady;
		this.Chan6TxFifoReady = this.HSSI_STAT1.Chan6TxFifoReady;
		this.HSSI_STAT1_Chan6RxDigitalResetTimeout = this.HSSI_STAT1.Chan6RxDigitalResetTimeout;
		this.Chan6RxDigitalResetTimeout = this.HSSI_STAT1.Chan6RxDigitalResetTimeout;
		this.HSSI_STAT1_Chan6TxDigitalResetTimeout = this.HSSI_STAT1.Chan6TxDigitalResetTimeout;
		this.Chan6TxDigitalResetTimeout = this.HSSI_STAT1.Chan6TxDigitalResetTimeout;
		this.HSSI_STAT1_Chan6RxDigitalResetStat = this.HSSI_STAT1.Chan6RxDigitalResetStat;
		this.Chan6RxDigitalResetStat = this.HSSI_STAT1.Chan6RxDigitalResetStat;
		this.HSSI_STAT1_Chan6RxAnalogResetStat = this.HSSI_STAT1.Chan6RxAnalogResetStat;
		this.Chan6RxAnalogResetStat = this.HSSI_STAT1.Chan6RxAnalogResetStat;
		this.HSSI_STAT1_Chan6TxDigitalResetStat = this.HSSI_STAT1.Chan6TxDigitalResetStat;
		this.Chan6TxDigitalResetStat = this.HSSI_STAT1.Chan6TxDigitalResetStat;
		this.HSSI_STAT1_Chan6TxAnalogResetStat = this.HSSI_STAT1.Chan6TxAnalogResetStat;
		this.Chan6TxAnalogResetStat = this.HSSI_STAT1.Chan6TxAnalogResetStat;
		this.HSSI_STAT1_Chan5RxReady = this.HSSI_STAT1.Chan5RxReady;
		this.Chan5RxReady = this.HSSI_STAT1.Chan5RxReady;
		this.HSSI_STAT1_Chan5TxReady = this.HSSI_STAT1.Chan5TxReady;
		this.Chan5TxReady = this.HSSI_STAT1.Chan5TxReady;
		this.HSSI_STAT1_Chan5RxIsLockedToRef = this.HSSI_STAT1.Chan5RxIsLockedToRef;
		this.Chan5RxIsLockedToRef = this.HSSI_STAT1.Chan5RxIsLockedToRef;
		this.HSSI_STAT1_Chan5RxIsLockedToData = this.HSSI_STAT1.Chan5RxIsLockedToData;
		this.Chan5RxIsLockedToData = this.HSSI_STAT1.Chan5RxIsLockedToData;
		this.HSSI_STAT1_Chan5RxCalBusy = this.HSSI_STAT1.Chan5RxCalBusy;
		this.Chan5RxCalBusy = this.HSSI_STAT1.Chan5RxCalBusy;
		this.HSSI_STAT1_Chan1TxCalBusy = this.HSSI_STAT1.Chan1TxCalBusy;
		this.HSSI_STAT1_Chan5RxTransferReady = this.HSSI_STAT1.Chan5RxTransferReady;
		this.Chan5RxTransferReady = this.HSSI_STAT1.Chan5RxTransferReady;
		this.HSSI_STAT1_Chan5TxTransferReady = this.HSSI_STAT1.Chan5TxTransferReady;
		this.Chan5TxTransferReady = this.HSSI_STAT1.Chan5TxTransferReady;
		this.HSSI_STAT1_Chan5RxFifoReady = this.HSSI_STAT1.Chan5RxFifoReady;
		this.Chan5RxFifoReady = this.HSSI_STAT1.Chan5RxFifoReady;
		this.HSSI_STAT1_Chan5TxFifoReady = this.HSSI_STAT1.Chan5TxFifoReady;
		this.Chan5TxFifoReady = this.HSSI_STAT1.Chan5TxFifoReady;
		this.HSSI_STAT1_Chan5RxDigitalResetTimeout = this.HSSI_STAT1.Chan5RxDigitalResetTimeout;
		this.Chan5RxDigitalResetTimeout = this.HSSI_STAT1.Chan5RxDigitalResetTimeout;
		this.HSSI_STAT1_Chan5TxDigitalResetTimeout = this.HSSI_STAT1.Chan5TxDigitalResetTimeout;
		this.Chan5TxDigitalResetTimeout = this.HSSI_STAT1.Chan5TxDigitalResetTimeout;
		this.HSSI_STAT1_Chan5RxDigitalResetStat = this.HSSI_STAT1.Chan5RxDigitalResetStat;
		this.Chan5RxDigitalResetStat = this.HSSI_STAT1.Chan5RxDigitalResetStat;
		this.HSSI_STAT1_Chan5RxAnalogResetStat = this.HSSI_STAT1.Chan5RxAnalogResetStat;
		this.Chan5RxAnalogResetStat = this.HSSI_STAT1.Chan5RxAnalogResetStat;
		this.HSSI_STAT1_Chan5TxDigitalResetStat = this.HSSI_STAT1.Chan5TxDigitalResetStat;
		this.Chan5TxDigitalResetStat = this.HSSI_STAT1.Chan5TxDigitalResetStat;
		this.HSSI_STAT1_Chan5TxAnalogResetStat = this.HSSI_STAT1.Chan5TxAnalogResetStat;
		this.Chan5TxAnalogResetStat = this.HSSI_STAT1.Chan5TxAnalogResetStat;
		this.HSSI_STAT1_Chan4RxReady = this.HSSI_STAT1.Chan4RxReady;
		this.Chan4RxReady = this.HSSI_STAT1.Chan4RxReady;
		this.HSSI_STAT1_Chan4TxReady = this.HSSI_STAT1.Chan4TxReady;
		this.Chan4TxReady = this.HSSI_STAT1.Chan4TxReady;
		this.HSSI_STAT1_Chan4RxIsLockedToRef = this.HSSI_STAT1.Chan4RxIsLockedToRef;
		this.Chan4RxIsLockedToRef = this.HSSI_STAT1.Chan4RxIsLockedToRef;
		this.HSSI_STAT1_Chan4RxIsLockedToData = this.HSSI_STAT1.Chan4RxIsLockedToData;
		this.Chan4RxIsLockedToData = this.HSSI_STAT1.Chan4RxIsLockedToData;
		this.HSSI_STAT1_Chan4RxCalBusy = this.HSSI_STAT1.Chan4RxCalBusy;
		this.Chan4RxCalBusy = this.HSSI_STAT1.Chan4RxCalBusy;
		this.HSSI_STAT1_Chan4TxCalBusy = this.HSSI_STAT1.Chan4TxCalBusy;
		this.Chan4TxCalBusy = this.HSSI_STAT1.Chan4TxCalBusy;
		this.HSSI_STAT1_Chan4RxTransferReady = this.HSSI_STAT1.Chan4RxTransferReady;
		this.Chan4RxTransferReady = this.HSSI_STAT1.Chan4RxTransferReady;
		this.HSSI_STAT1_Chan4TxTransferReady = this.HSSI_STAT1.Chan4TxTransferReady;
		this.Chan4TxTransferReady = this.HSSI_STAT1.Chan4TxTransferReady;
		this.HSSI_STAT1_Chan4RxFifoReady = this.HSSI_STAT1.Chan4RxFifoReady;
		this.Chan4RxFifoReady = this.HSSI_STAT1.Chan4RxFifoReady;
		this.HSSI_STAT1_Chan4TxFifoReady = this.HSSI_STAT1.Chan4TxFifoReady;
		this.Chan4TxFifoReady = this.HSSI_STAT1.Chan4TxFifoReady;
		this.HSSI_STAT1_Chan4RxDigitalResetTimeout = this.HSSI_STAT1.Chan4RxDigitalResetTimeout;
		this.Chan4RxDigitalResetTimeout = this.HSSI_STAT1.Chan4RxDigitalResetTimeout;
		this.HSSI_STAT1_Chan4TxDigitalResetTimeout = this.HSSI_STAT1.Chan4TxDigitalResetTimeout;
		this.Chan4TxDigitalResetTimeout = this.HSSI_STAT1.Chan4TxDigitalResetTimeout;
		this.HSSI_STAT1_Chan4RxDigitalResetStat = this.HSSI_STAT1.Chan4RxDigitalResetStat;
		this.Chan4RxDigitalResetStat = this.HSSI_STAT1.Chan4RxDigitalResetStat;
		this.HSSI_STAT1_Chan4RxAnalogResetStat = this.HSSI_STAT1.Chan4RxAnalogResetStat;
		this.Chan4RxAnalogResetStat = this.HSSI_STAT1.Chan4RxAnalogResetStat;
		this.HSSI_STAT1_Chan4TxDigitalResetStat = this.HSSI_STAT1.Chan4TxDigitalResetStat;
		this.Chan4TxDigitalResetStat = this.HSSI_STAT1.Chan4TxDigitalResetStat;
		this.HSSI_STAT1_Chan4TxAnalogResetStat = this.HSSI_STAT1.Chan4TxAnalogResetStat;
		this.Chan4TxAnalogResetStat = this.HSSI_STAT1.Chan4TxAnalogResetStat;
      this.HSSI_RCFG_CMD0 = ral_reg_hssi_ss_csr_HSSI_RCFG_CMD0::type_id::create("HSSI_RCFG_CMD0",,get_full_name());
      this.HSSI_RCFG_CMD0.configure(this, null, "");
      this.HSSI_RCFG_CMD0.build();
      this.default_map.add_reg(this.HSSI_RCFG_CMD0, `UVM_REG_ADDR_WIDTH'h28, "RW", 0);
		this.HSSI_RCFG_CMD0_Reserved = this.HSSI_RCFG_CMD0.Reserved;
		this.HSSI_RCFG_CMD0_XcvrRcfgAddr = this.HSSI_RCFG_CMD0.XcvrRcfgAddr;
		this.XcvrRcfgAddr = this.HSSI_RCFG_CMD0.XcvrRcfgAddr;
		this.HSSI_RCFG_CMD0_Reserved_1 = this.HSSI_RCFG_CMD0.Reserved_1;
		this.Reserved_1 = this.HSSI_RCFG_CMD0.Reserved_1;
		this.HSSI_RCFG_CMD0_XcvrRcfgAck = this.HSSI_RCFG_CMD0.XcvrRcfgAck;
		this.XcvrRcfgAck = this.HSSI_RCFG_CMD0.XcvrRcfgAck;
		this.HSSI_RCFG_CMD0_XcvrRcfgCmdStatus = this.HSSI_RCFG_CMD0.XcvrRcfgCmdStatus;
		this.XcvrRcfgCmdStatus = this.HSSI_RCFG_CMD0.XcvrRcfgCmdStatus;
      this.HSSI_RCFG_DATA0 = ral_reg_hssi_ss_csr_HSSI_RCFG_DATA0::type_id::create("HSSI_RCFG_DATA0",,get_full_name());
      this.HSSI_RCFG_DATA0.configure(this, null, "");
      this.HSSI_RCFG_DATA0.build();
      this.default_map.add_reg(this.HSSI_RCFG_DATA0, `UVM_REG_ADDR_WIDTH'h30, "RW", 0);
		this.HSSI_RCFG_DATA0_XcvrRcfgWrData = this.HSSI_RCFG_DATA0.XcvrRcfgWrData;
		this.XcvrRcfgWrData = this.HSSI_RCFG_DATA0.XcvrRcfgWrData;
		this.HSSI_RCFG_DATA0_XcvrRcfgRdData = this.HSSI_RCFG_DATA0.XcvrRcfgRdData;
		this.XcvrRcfgRdData = this.HSSI_RCFG_DATA0.XcvrRcfgRdData;
      this.HSSI_SCRATCHPAD = ral_reg_hssi_ss_csr_HSSI_SCRATCHPAD::type_id::create("HSSI_SCRATCHPAD",,get_full_name());
      this.HSSI_SCRATCHPAD.configure(this, null, "");
      this.HSSI_SCRATCHPAD.build();
      this.default_map.add_reg(this.HSSI_SCRATCHPAD, `UVM_REG_ADDR_WIDTH'h38, "RW", 0);
		this.HSSI_SCRATCHPAD_Scrathpad = this.HSSI_SCRATCHPAD.Scrathpad;
		this.Scrathpad = this.HSSI_SCRATCHPAD.Scrathpad;
   endfunction : build

	`uvm_object_utils(ral_block_hssi_ss_csr)

endclass : ral_block_hssi_ss_csr



`endif
